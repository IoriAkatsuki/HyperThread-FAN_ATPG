module TC01 (
test_siA,
test_seA,
test_soA,
CKA,
g18A,
g27A,
g109A,
g741A,
g742A,
g743A,
g744A,
g872A,
g873A,
g877A,
g881A,
g1712A,
g1960A,
g1961A,
g1696A,
g750A,
g85A,
g42A,
g1700A,
g102A,
g104A,
g101A,
g29A,
g28A,
g103A,
g83A,
g23A,
g87A,
g922A,
g892A,
g84A,
g919A,
g1182A,
g925A,
g48A,
g895A,
g889A,
g1185A,
g41A,
g43A,
g99A,
g1173A,
g1203A,
g1188A,
g1197A,
g46A,
g31A,
g45A,
g92A,
g89A,
g898A,
g91A,
g93A,
g913A,
g82A,
g88A,
g1194A,
g47A,
g96A,
g910A,
g95A,
g904A,
g1176A,
g901A,
g44A,
g916A,
g100A,
g886A,
g30A,
g86A,
g1170A,
g1200A,
g1191A,
g907A,
g90A,
g94A,
g1179A,
g2355A,
g2601A,
g2602A,
g2603A,
g2604A,
g2605A,
g2606A,
g2607A,
g2608A,
g2609A,
g2610A,
g2611A,
g2612A,
g2648A,
g2986A,
g3007A,
g3069A,
g4172A,
g4173A,
g4174A,
g4175A,
g4176A,
g4177A,
g4178A,
g4179A,
g4180A,
g4181A,
g4887A,
g4888A,
g5101A,
g5105A,
g5658A,
g5659A,
g5816A,
g6920A,
g6926A,
g6932A,
g6942A,
g6949A,
g6955A,
g7744A,
g8061A,
g8062A,
g8271A,
g8313A,
g8316A,
g8318A,
g8323A,
g8328A,
g8331A,
g8335A,
g8340A,
g8347A,
g8349A,
g8352A,
g8561A,
g8562A,
g8563A,
g8564A,
g8565A,
g8566A,
g8976A,
g8977A,
g8978A,
g8979A,
g8980A,
g8981A,
g8982A,
g8983A,
g8984A,
g8985A,
g8986A,
g9451A,
g9961A,
g10377A,
g10379A,
g10455A,
g10457A,
g10459A,
g10461A,
g10463A,
g10465A,
g10628A,
g10801A,
g11163A,
g11206A,
g11489A,
g6842A,
g4171A,
g6267A,
g6257A,
g1957A,
g6282A,
g6284A,
g6281A,
g6253A,
g6285A,
g6283A,
g6265A,
g3327A,
g6269A,
g4204A,
g4193A,
g6266A,
g4203A,
g4212A,
g4196A,
g6263A,
g4194A,
g4192A,
g4213A,
g6256A,
g6258A,
g6279A,
g4209A,
g4208A,
g4214A,
g4206A,
g6261A,
g6255A,
g6260A,
g6274A,
g6271A,
g4195A,
g6273A,
g6275A,
g4201A,
g6264A,
g6270A,
g4216A,
g6262A,
g6278A,
g4200A,
g6277A,
g4198A,
g4210A,
g4197A,
g6259A,
g4202A,
g6280A,
g4191A,
g6254A,
g6268A,
g4205A,
g4207A,
g4215A,
g4199A,
g6272A,
g6276A,
g4211A,
test_siB,
test_seB,
test_soB,
CKB,
g18B,
g27B,
g109B,
g741B,
g742B,
g743B,
g744B,
g872B,
g873B,
g877B,
g881B,
g1712B,
g1960B,
g1961B,
g1696B,
g750B,
g85B,
g42B,
g1700B,
g102B,
g104B,
g101B,
g29B,
g28B,
g103B,
g83B,
g23B,
g87B,
g922B,
g892B,
g84B,
g919B,
g1182B,
g925B,
g48B,
g895B,
g889B,
g1185B,
g41B,
g43B,
g99B,
g1173B,
g1203B,
g1188B,
g1197B,
g46B,
g31B,
g45B,
g92B,
g89B,
g898B,
g91B,
g93B,
g913B,
g82B,
g88B,
g1194B,
g47B,
g96B,
g910B,
g95B,
g904B,
g1176B,
g901B,
g44B,
g916B,
g100B,
g886B,
g30B,
g86B,
g1170B,
g1200B,
g1191B,
g907B,
g90B,
g94B,
g1179B,
g2355B,
g2601B,
g2602B,
g2603B,
g2604B,
g2605B,
g2606B,
g2607B,
g2608B,
g2609B,
g2610B,
g2611B,
g2612B,
g2648B,
g2986B,
g3007B,
g3069B,
g4172B,
g4173B,
g4174B,
g4175B,
g4176B,
g4177B,
g4178B,
g4179B,
g4180B,
g4181B,
g4887B,
g4888B,
g5101B,
g5105B,
g5658B,
g5659B,
g5816B,
g6920B,
g6926B,
g6932B,
g6942B,
g6949B,
g6955B,
g7744B,
g8061B,
g8062B,
g8271B,
g8313B,
g8316B,
g8318B,
g8323B,
g8328B,
g8331B,
g8335B,
g8340B,
g8347B,
g8349B,
g8352B,
g8561B,
g8562B,
g8563B,
g8564B,
g8565B,
g8566B,
g8976B,
g8977B,
g8978B,
g8979B,
g8980B,
g8981B,
g8982B,
g8983B,
g8984B,
g8985B,
g8986B,
g9451B,
g9961B,
g10377B,
g10379B,
g10455B,
g10457B,
g10459B,
g10461B,
g10463B,
g10465B,
g10628B,
g10801B,
g11163B,
g11206B,
g11489B,
g6842B,
g4171B,
g6267B,
g6257B,
g1957B,
g6282B,
g6284B,
g6281B,
g6253B,
g6285B,
g6283B,
g6265B,
g3327B,
g6269B,
g4204B,
g4193B,
g6266B,
g4203B,
g4212B,
g4196B,
g6263B,
g4194B,
g4192B,
g4213B,
g6256B,
g6258B,
g6279B,
g4209B,
g4208B,
g4214B,
g4206B,
g6261B,
g6255B,
g6260B,
g6274B,
g6271B,
g4195B,
g6273B,
g6275B,
g4201B,
g6264B,
g6270B,
g4216B,
g6262B,
g6278B,
g4200B,
g6277B,
g4198B,
g4210B,
g4197B,
g6259B,
g4202B,
g6280B,
g4191B,
g6254B,
g6268B,
g4205B,
g4207B,
g4215B,
g4199B,
g6272B,
g6276B,
g4211B,
test_siC,
test_seC,
test_soC,
CKC,
g18C,
g27C,
g109C,
g741C,
g742C,
g743C,
g744C,
g872C,
g873C,
g877C,
g881C,
g1712C,
g1960C,
g1961C,
g1696C,
g750C,
g85C,
g42C,
g1700C,
g102C,
g104C,
g101C,
g29C,
g28C,
g103C,
g83C,
g23C,
g87C,
g922C,
g892C,
g84C,
g919C,
g1182C,
g925C,
g48C,
g895C,
g889C,
g1185C,
g41C,
g43C,
g99C,
g1173C,
g1203C,
g1188C,
g1197C,
g46C,
g31C,
g45C,
g92C,
g89C,
g898C,
g91C,
g93C,
g913C,
g82C,
g88C,
g1194C,
g47C,
g96C,
g910C,
g95C,
g904C,
g1176C,
g901C,
g44C,
g916C,
g100C,
g886C,
g30C,
g86C,
g1170C,
g1200C,
g1191C,
g907C,
g90C,
g94C,
g1179C,
g2355C,
g2601C,
g2602C,
g2603C,
g2604C,
g2605C,
g2606C,
g2607C,
g2608C,
g2609C,
g2610C,
g2611C,
g2612C,
g2648C,
g2986C,
g3007C,
g3069C,
g4172C,
g4173C,
g4174C,
g4175C,
g4176C,
g4177C,
g4178C,
g4179C,
g4180C,
g4181C,
g4887C,
g4888C,
g5101C,
g5105C,
g5658C,
g5659C,
g5816C,
g6920C,
g6926C,
g6932C,
g6942C,
g6949C,
g6955C,
g7744C,
g8061C,
g8062C,
g8271C,
g8313C,
g8316C,
g8318C,
g8323C,
g8328C,
g8331C,
g8335C,
g8340C,
g8347C,
g8349C,
g8352C,
g8561C,
g8562C,
g8563C,
g8564C,
g8565C,
g8566C,
g8976C,
g8977C,
g8978C,
g8979C,
g8980C,
g8981C,
g8982C,
g8983C,
g8984C,
g8985C,
g8986C,
g9451C,
g9961C,
g10377C,
g10379C,
g10455C,
g10457C,
g10459C,
g10461C,
g10463C,
g10465C,
g10628C,
g10801C,
g11163C,
g11206C,
g11489C,
g6842C,
g4171C,
g6267C,
g6257C,
g1957C,
g6282C,
g6284C,
g6281C,
g6253C,
g6285C,
g6283C,
g6265C,
g3327C,
g6269C,
g4204C,
g4193C,
g6266C,
g4203C,
g4212C,
g4196C,
g6263C,
g4194C,
g4192C,
g4213C,
g6256C,
g6258C,
g6279C,
g4209C,
g4208C,
g4214C,
g4206C,
g6261C,
g6255C,
g6260C,
g6274C,
g6271C,
g4195C,
g6273C,
g6275C,
g4201C,
g6264C,
g6270C,
g4216C,
g6262C,
g6278C,
g4200C,
g6277C,
g4198C,
g4210C,
g4197C,
g6259C,
g4202C,
g6280C,
g4191C,
g6254C,
g6268C,
g4205C,
g4207C,
g4215C,
g4199C,
g6272C,
g6276C,
g4211C);
input CKA;
input test_siA;
input test_seA;
output test_soA;
input g18A;
input g27A;
input g109A;
input g741A;
input g742A;
input g743A;
input g744A;
input g872A;
input g873A;
input g877A;
input g881A;
input g1712A;
input g1960A;
input g1961A;
input g1696A;
input g750A;
input g85A;
input g42A;
input g1700A;
input g102A;
input g104A;
input g101A;
input g29A;
input g28A;
input g103A;
input g83A;
input g23A;
input g87A;
input g922A;
input g892A;
input g84A;
input g919A;
input g1182A;
input g925A;
input g48A;
input g895A;
input g889A;
input g1185A;
input g41A;
input g43A;
input g99A;
input g1173A;
input g1203A;
input g1188A;
input g1197A;
input g46A;
input g31A;
input g45A;
input g92A;
input g89A;
input g898A;
input g91A;
input g93A;
input g913A;
input g82A;
input g88A;
input g1194A;
input g47A;
input g96A;
input g910A;
input g95A;
input g904A;
input g1176A;
input g901A;
input g44A;
input g916A;
input g100A;
input g886A;
input g30A;
input g86A;
input g1170A;
input g1200A;
input g1191A;
input g907A;
input g90A;
input g94A;
input g1179A;
output g2355A;
output g2601A;
output g2602A;
output g2603A;
output g2604A;
output g2605A;
output g2606A;
output g2607A;
output g2608A;
output g2609A;
output g2610A;
output g2611A;
output g2612A;
output g2648A;
output g2986A;
output g3007A;
output g3069A;
output g4172A;
output g4173A;
output g4174A;
output g4175A;
output g4176A;
output g4177A;
output g4178A;
output g4179A;
output g4180A;
output g4181A;
output g4887A;
output g4888A;
output g5101A;
output g5105A;
output g5658A;
output g5659A;
output g5816A;
output g6920A;
output g6926A;
output g6932A;
output g6942A;
output g6949A;
output g6955A;
output g7744A;
output g8061A;
output g8062A;
output g8271A;
output g8313A;
output g8316A;
output g8318A;
output g8323A;
output g8328A;
output g8331A;
output g8335A;
output g8340A;
output g8347A;
output g8349A;
output g8352A;
output g8561A;
output g8562A;
output g8563A;
output g8564A;
output g8565A;
output g8566A;
output g8976A;
output g8977A;
output g8978A;
output g8979A;
output g8980A;
output g8981A;
output g8982A;
output g8983A;
output g8984A;
output g8985A;
output g8986A;
output g9451A;
output g9961A;
output g10377A;
output g10379A;
output g10455A;
output g10457A;
output g10459A;
output g10461A;
output g10463A;
output g10465A;
output g10628A;
output g10801A;
output g11163A;
output g11206A;
output g11489A;
output g6842A;
output g4171A;
output g6267A;
output g6257A;
output g1957A;
output g6282A;
output g6284A;
output g6281A;
output g6253A;
output g6285A;
output g6283A;
output g6265A;
output g3327A;
output g6269A;
output g4204A;
output g4193A;
output g6266A;
output g4203A;
output g4212A;
output g4196A;
output g6263A;
output g4194A;
output g4192A;
output g4213A;
output g6256A;
output g6258A;
output g6279A;
output g4209A;
output g4208A;
output g4214A;
output g4206A;
output g6261A;
output g6255A;
output g6260A;
output g6274A;
output g6271A;
output g4195A;
output g6273A;
output g6275A;
output g4201A;
output g6264A;
output g6270A;
output g4216A;
output g6262A;
output g6278A;
output g4200A;
output g6277A;
output g4198A;
output g4210A;
output g4197A;
output g6259A;
output g4202A;
output g6280A;
output g4191A;
output g6254A;
output g6268A;
output g4205A;
output g4207A;
output g4215A;
output g4199A;
output g6272A;
output g6276A;
output g4211A;
input CKB;
input test_siB;
input test_seB;
output test_soB;
input g18B;
input g27B;
input g109B;
input g741B;
input g742B;
input g743B;
input g744B;
input g872B;
input g873B;
input g877B;
input g881B;
input g1712B;
input g1960B;
input g1961B;
input g1696B;
input g750B;
input g85B;
input g42B;
input g1700B;
input g102B;
input g104B;
input g101B;
input g29B;
input g28B;
input g103B;
input g83B;
input g23B;
input g87B;
input g922B;
input g892B;
input g84B;
input g919B;
input g1182B;
input g925B;
input g48B;
input g895B;
input g889B;
input g1185B;
input g41B;
input g43B;
input g99B;
input g1173B;
input g1203B;
input g1188B;
input g1197B;
input g46B;
input g31B;
input g45B;
input g92B;
input g89B;
input g898B;
input g91B;
input g93B;
input g913B;
input g82B;
input g88B;
input g1194B;
input g47B;
input g96B;
input g910B;
input g95B;
input g904B;
input g1176B;
input g901B;
input g44B;
input g916B;
input g100B;
input g886B;
input g30B;
input g86B;
input g1170B;
input g1200B;
input g1191B;
input g907B;
input g90B;
input g94B;
input g1179B;
output g2355B;
output g2601B;
output g2602B;
output g2603B;
output g2604B;
output g2605B;
output g2606B;
output g2607B;
output g2608B;
output g2609B;
output g2610B;
output g2611B;
output g2612B;
output g2648B;
output g2986B;
output g3007B;
output g3069B;
output g4172B;
output g4173B;
output g4174B;
output g4175B;
output g4176B;
output g4177B;
output g4178B;
output g4179B;
output g4180B;
output g4181B;
output g4887B;
output g4888B;
output g5101B;
output g5105B;
output g5658B;
output g5659B;
output g5816B;
output g6920B;
output g6926B;
output g6932B;
output g6942B;
output g6949B;
output g6955B;
output g7744B;
output g8061B;
output g8062B;
output g8271B;
output g8313B;
output g8316B;
output g8318B;
output g8323B;
output g8328B;
output g8331B;
output g8335B;
output g8340B;
output g8347B;
output g8349B;
output g8352B;
output g8561B;
output g8562B;
output g8563B;
output g8564B;
output g8565B;
output g8566B;
output g8976B;
output g8977B;
output g8978B;
output g8979B;
output g8980B;
output g8981B;
output g8982B;
output g8983B;
output g8984B;
output g8985B;
output g8986B;
output g9451B;
output g9961B;
output g10377B;
output g10379B;
output g10455B;
output g10457B;
output g10459B;
output g10461B;
output g10463B;
output g10465B;
output g10628B;
output g10801B;
output g11163B;
output g11206B;
output g11489B;
output g6842B;
output g4171B;
output g6267B;
output g6257B;
output g1957B;
output g6282B;
output g6284B;
output g6281B;
output g6253B;
output g6285B;
output g6283B;
output g6265B;
output g3327B;
output g6269B;
output g4204B;
output g4193B;
output g6266B;
output g4203B;
output g4212B;
output g4196B;
output g6263B;
output g4194B;
output g4192B;
output g4213B;
output g6256B;
output g6258B;
output g6279B;
output g4209B;
output g4208B;
output g4214B;
output g4206B;
output g6261B;
output g6255B;
output g6260B;
output g6274B;
output g6271B;
output g4195B;
output g6273B;
output g6275B;
output g4201B;
output g6264B;
output g6270B;
output g4216B;
output g6262B;
output g6278B;
output g4200B;
output g6277B;
output g4198B;
output g4210B;
output g4197B;
output g6259B;
output g4202B;
output g6280B;
output g4191B;
output g6254B;
output g6268B;
output g4205B;
output g4207B;
output g4215B;
output g4199B;
output g6272B;
output g6276B;
output g4211B;
input CKC;
input test_siC;
input test_seC;
output test_soC;
input g18C;
input g27C;
input g109C;
input g741C;
input g742C;
input g743C;
input g744C;
input g872C;
input g873C;
input g877C;
input g881C;
input g1712C;
input g1960C;
input g1961C;
input g1696C;
input g750C;
input g85C;
input g42C;
input g1700C;
input g102C;
input g104C;
input g101C;
input g29C;
input g28C;
input g103C;
input g83C;
input g23C;
input g87C;
input g922C;
input g892C;
input g84C;
input g919C;
input g1182C;
input g925C;
input g48C;
input g895C;
input g889C;
input g1185C;
input g41C;
input g43C;
input g99C;
input g1173C;
input g1203C;
input g1188C;
input g1197C;
input g46C;
input g31C;
input g45C;
input g92C;
input g89C;
input g898C;
input g91C;
input g93C;
input g913C;
input g82C;
input g88C;
input g1194C;
input g47C;
input g96C;
input g910C;
input g95C;
input g904C;
input g1176C;
input g901C;
input g44C;
input g916C;
input g100C;
input g886C;
input g30C;
input g86C;
input g1170C;
input g1200C;
input g1191C;
input g907C;
input g90C;
input g94C;
input g1179C;
output g2355C;
output g2601C;
output g2602C;
output g2603C;
output g2604C;
output g2605C;
output g2606C;
output g2607C;
output g2608C;
output g2609C;
output g2610C;
output g2611C;
output g2612C;
output g2648C;
output g2986C;
output g3007C;
output g3069C;
output g4172C;
output g4173C;
output g4174C;
output g4175C;
output g4176C;
output g4177C;
output g4178C;
output g4179C;
output g4180C;
output g4181C;
output g4887C;
output g4888C;
output g5101C;
output g5105C;
output g5658C;
output g5659C;
output g5816C;
output g6920C;
output g6926C;
output g6932C;
output g6942C;
output g6949C;
output g6955C;
output g7744C;
output g8061C;
output g8062C;
output g8271C;
output g8313C;
output g8316C;
output g8318C;
output g8323C;
output g8328C;
output g8331C;
output g8335C;
output g8340C;
output g8347C;
output g8349C;
output g8352C;
output g8561C;
output g8562C;
output g8563C;
output g8564C;
output g8565C;
output g8566C;
output g8976C;
output g8977C;
output g8978C;
output g8979C;
output g8980C;
output g8981C;
output g8982C;
output g8983C;
output g8984C;
output g8985C;
output g8986C;
output g9451C;
output g9961C;
output g10377C;
output g10379C;
output g10455C;
output g10457C;
output g10459C;
output g10461C;
output g10463C;
output g10465C;
output g10628C;
output g10801C;
output g11163C;
output g11206C;
output g11489C;
output g6842C;
output g4171C;
output g6267C;
output g6257C;
output g1957C;
output g6282C;
output g6284C;
output g6281C;
output g6253C;
output g6285C;
output g6283C;
output g6265C;
output g3327C;
output g6269C;
output g4204C;
output g4193C;
output g6266C;
output g4203C;
output g4212C;
output g4196C;
output g6263C;
output g4194C;
output g4192C;
output g4213C;
output g6256C;
output g6258C;
output g6279C;
output g4209C;
output g4208C;
output g4214C;
output g4206C;
output g6261C;
output g6255C;
output g6260C;
output g6274C;
output g6271C;
output g4195C;
output g6273C;
output g6275C;
output g4201C;
output g6264C;
output g6270C;
output g4216C;
output g6262C;
output g6278C;
output g4200C;
output g6277C;
output g4198C;
output g4210C;
output g4197C;
output g6259C;
output g4202C;
output g6280C;
output g4191C;
output g6254C;
output g6268C;
output g4205C;
output g4207C;
output g4215C;
output g4199C;
output g6272C;
output g6276C;
output g4211C;

   // Internal wires
wire FE_OFN370_g4525A;
wire FE_OFN369_g4525A;
wire FE_OFN368_g4525A;
wire FE_OFN367_g3521A;
wire FE_OFN366_g3521A;
wire FE_OFN365_g5361A;
wire FE_OFN364_g3015A;
wire FE_OFN363_I5565A;
wire FE_OFN362_g4525A;
wire FE_OFN360_g4525A;
wire FE_OFN359_g18A;
wire FE_OFN358_g3521A;
wire FE_OFN357_g3521A;
wire FE_OFN356_g5361A;
wire FE_OFN354_g5361A;
wire FE_OFN353_g5117A;
wire FE_OFN352_g109A;
wire FE_OFN351_g3913A;
wire FE_OFN350_g3121A;
wire FE_OFN349_I6424A;
wire FE_OFN348_g3015A;
wire FE_OFN347_g3914A;
wire FE_OFN346_g4381A;
wire FE_OFN345_g3015A;
wire FE_OFN344_g3586A;
wire FE_OFN343_I5565A;
wire FE_OFN340_I5565A;
wire FE_OFN339_g4525A;
wire FE_OFN337_g4525A;
wire FE_OFN336_g1690A;
wire FE_OFN335_g4737A;
wire FE_OFN334_g7045A;
wire FE_OFN333_g4294A;
wire FE_OFN332_g8748A;
wire FE_OFN331_g8696A;
wire FE_OFN330_g7638A;
wire FE_OFN329_g8763A;
wire FE_OFN328_g8709A;
wire FE_OFN325_g18A;
wire FE_OFN324_g18A;
wire FE_OFN322_g4449A;
wire FE_OFN321_g5261A;
wire FE_OFN320_g5361A;
wire FE_OFN319_g5361A;
wire FE_OFN318_g5361A;
wire FE_OFN316_g5361A;
wire FE_OFN315_g5117A;
wire FE_OFN312_g5117A;
wire FE_OFN310_g4336A;
wire FE_OFN308_I6424A;
wire FE_OFN307_g4010A;
wire FE_OFN306_g5128A;
wire FE_OFN305_g5151A;
wire FE_OFN304_g5151A;
wire FE_OFN303_g4678A;
wire FE_OFN302_g3913A;
wire FE_OFN300_g4002A;
wire FE_OFN299_g4457A;
wire FE_OFN298_g3015A;
wire FE_OFN297_g3015A;
wire FE_OFN296_g3914A;
wire FE_OFN294_g3914A;
wire FE_OFN293_g3015A;
wire FE_OFN292_g3015A;
wire FE_OFN291_g4880A;
wire FE_OFN290_g4880A;
wire FE_OFN289_g4679A;
wire FE_OFN288_g4263A;
wire FE_OFN287_g3586A;
wire FE_OFN284_g3586A;
wire FE_OFN283_I8869A;
wire FE_OFN282_g6165A;
wire FE_OFN281_g2216A;
wire FE_OFN280_g9536A;
wire FE_OFN279_g11157A;
wire FE_OFN278_g10927A;
wire FE_OFN277_g48A;
wire FE_OFN276_g48A;
wire FE_OFN275_g48A;
wire FE_OFN273_g85A;
wire FE_OFN271_g85A;
wire FE_OFN269_g109A;
wire FE_OFN267_g109A;
wire FE_OFN266_g18A;
wire FE_OFN260_g18A;
wire FE_OFN254_g461A;
wire FE_OFN253_g1786A;
wire FE_OFN252_g1791A;
wire FE_OFN251_g1801A;
wire FE_OFN250_g471A;
wire FE_OFN248_g466A;
wire FE_OFN247_g1771A;
wire FE_OFN245_g1690A;
wire FE_OFN241_g1690A;
wire FE_OFN240_g1110A;
wire FE_OFN239_g1796A;
wire FE_OFN238_g1781A;
wire FE_OFN237_g1806A;
wire FE_OFN236_g1776A;
wire FE_OFN235_g2024A;
wire FE_OFN234_g2024A;
wire FE_OFN233_I5565A;
wire FE_OFN230_I5565A;
wire FE_OFN229_g3880A;
wire FE_OFN227_g3880A;
wire FE_OFN226_g3880A;
wire FE_OFN225_g2276A;
wire FE_OFN224_g2276A;
wire FE_OFN223_g4401A;
wire FE_OFN221_g3440A;
wire FE_OFN219_g5557A;
wire FE_OFN218_g5557A;
wire FE_OFN217_g5013A;
wire FE_OFN213_g6003A;
wire FE_OFN211_g7246A;
wire FE_OFN210_g7246A;
wire FE_OFN209_g6863A;
wire FE_OFN207_g6863A;
wire FE_OFN206_g6863A;
wire FE_OFN204_g3664A;
wire FE_OFN200_g4921A;
wire FE_OFN199_g7697A;
wire FE_OFN198_g7697A;
wire FE_OFN196_g7697A;
wire FE_OFN195_g6488A;
wire FE_OFN192_g6488A;
wire FE_OFN191_g6488A;
wire FE_OFN189_g7638A;
wire FE_OFN187_g7638A;
wire FE_OFN184_I7048A;
wire FE_OFN180_g5354A;
wire FE_OFN179_g5354A;
wire FE_OFN178_g5354A;
wire FE_OFN177_g5919A;
wire FE_OFN176_g5151A;
wire FE_OFN168_g5361A;
wire FE_OFN166_g5361A;
wire FE_OFN164_g5361A;
wire FE_OFN161_g5361A;
wire FE_OFN160_I6424A;
wire FE_OFN155_g3121A;
wire FE_OFN154_g4640A;
wire FE_OFN153_g4640A;
wire FE_OFN147_g4682A;
wire FE_OFN146_g4682A;
wire FE_OFN144_g4682A;
wire FE_OFN142_g4682A;
wire FE_OFN141_g3829A;
wire FE_OFN137_g3829A;
wire FE_OFN136_g3863A;
wire FE_OFN134_g3863A;
wire FE_OFN133_g3015A;
wire FE_OFN132_g3015A;
wire FE_OFN131_g3015A;
wire FE_OFN119_g3015A;
wire FE_OFN118_g4807A;
wire FE_OFN117_g4807A;
wire FE_OFN116_g4807A;
wire FE_OFN115_g4807A;
wire FE_OFN113_g3914A;
wire FE_OFN111_g3914A;
wire FE_OFN110_g3586A;
wire FE_OFN103_g3586A;
wire FE_OFN102_g3586A;
wire FE_OFN100_g4421A;
wire FE_OFN99_g4421A;
wire FE_OFN97_I8869A;
wire FE_OFN96_g2169A;
wire FE_OFN95_g2216A;
wire FE_OFN93_g2216A;
wire FE_OFN92_g2216A;
wire FE_OFN91_g2172A;
wire FE_OFN90_I11360A;
wire FE_OFN89_I11360A;
wire FE_OFN88_g2178A;
wire FE_OFN87_g2176A;
wire FE_OFN86_g2176A;
wire FE_OFN85_g2176A;
wire FE_OFN84_g2176A;
wire FE_OFN83_g2176A;
wire FE_OFN82_g2176A;
wire FE_OFN81_g2176A;
wire FE_OFN80_g2175A;
wire FE_OFN79_g8700A;
wire FE_OFN76_g8700A;
wire FE_OFN73_g8858A;
wire FE_OFN72_g9292A;
wire FE_OFN71_g9292A;
wire FE_OFN70_g9490A;
wire FE_OFN69_g9392A;
wire FE_OFN68_g9392A;
wire FE_OFN67_g9367A;
wire FE_OFN64_g9536A;
wire FE_OFN63_g9474A;
wire FE_OFN62_g9274A;
wire FE_OFN61_g9624A;
wire FE_OFN60_g9624A;
wire FE_OFN59_g9432A;
wire FE_OFN57_g9432A;
wire FE_OFN56_g9052A;
wire FE_OFN54_g9052A;
wire FE_OFN53_g9173A;
wire FE_OFN52_g9173A;
wire FE_OFN51_g9111A;
wire FE_OFN50_g9030A;
wire FE_OFN49_g9030A;
wire FE_OFN48_g9151A;
wire FE_OFN47_g9151A;
wire FE_OFN46_g9125A;
wire FE_OFN45_g9125A;
wire FE_OFN44_g9125A;
wire FE_OFN42_g9205A;
wire FE_OFN40_g9240A;
wire FE_OFN39_g9223A;
wire FE_OFN35_g9785A;
wire FE_OFN34_g9785A;
wire FE_OFN33_g9454A;
wire FE_OFN32_g9454A;
wire FE_OFN27_g11519A;
wire FE_OFN21_g10702A;
wire FE_OFN20_g10702A;
wire FE_OFN18_g10702A;
wire FE_OFN17_g10702A;
wire FE_OFN15_g10702A;
wire FE_OFN14_g10702A;
wire FE_OFN13_g10702A;
wire FE_OFN10_g10702A;
wire FE_OFN9_g10702A;
wire FE_OFN8_g10702A;
wire FE_OFN7_g10702A;
wire FE_OFN4_g10950A;
wire FE_OFN3_g10950A;
wire FE_OFN0_g10950A;
wire g4500A;
wire g5529A;
wire g9968A;
wire g4682A;
wire g1707A;
wire g2299A;
wire g9291A;
wire g2807A;
wire I7048A;
wire g4130A;
wire g5024A;
wire g4338A;
wire g11596A;
wire g8147A;
wire g6551A;
wire g10865A;
wire g650A;
wire g1981A;
wire g8054A;
wire g3982A;
wire g9974A;
wire g1216A;
wire g546A;
wire g798A;
wire g3629A;
wire g7709A;
wire g8465A;
wire g8617A;
wire g4940A;
wire g4640A;
wire g135A;
wire g2078A;
wire g4565A;
wire g1918A;
wire g2340A;
wire g7684A;
wire g11519A;
wire g5935A;
wire g3800A;
wire g4736A;
wire g6941A;
wire g201A;
wire g2435A;
wire g4010A;
wire g1371A;
wire g2082A;
wire g4811A;
wire g5519A;
wire g49A;
wire g560A;
wire g6481A;
wire g6215A;
wire g10563A;
wire g10668A;
wire g70A;
wire g5013A;
wire g11221A;
wire g9508A;
wire g5212A;
wire g6529A;
wire g8709A;
wire g115A;
wire g2214A;
wire g5008A;
wire g3829A;
wire g9995A;
wire g10707A;
wire g3435A;
wire I7847A;
wire g5576A;
wire I13400A;
wire I5002A;
wire g10013A;
wire g10385A;
wire g9432A;
wire g3753A;
wire g4566A;
wire g254A;
wire I14326A;
wire g4722A;
wire g3348A;
wire g9696A;
wire g10408A;
wire I15968A;
wire g756A;
wire g818A;
wire g10937A;
wire g11060A;
wire g7242A;
wire g10336A;
wire I15855A;
wire g5229A;
wire g8940A;
wire g259A;
wire g10584A;
wire g10679A;
wire g4560A;
wire g10855A;
wire g369A;
wire g1968A;
wire I15503A;
wire g7996A;
wire g8110A;
wire g186A;
wire g2556A;
wire g3586A;
wire g10496A;
wire g3399A;
wire I7817A;
wire g158A;
wire g2222A;
wire g6907A;
wire g8226A;
wire I13373A;
wire g5405A;
wire I9880A;
wire g6155A;
wire g7246A;
wire g6638A;
wire g11647A;
wire g2744A;
wire g4094A;
wire g32A;
wire g3374A;
wire g4567A;
wire g8814A;
wire I14312A;
wire g10950A;
wire g9490A;
wire g11111A;
wire g4776A;
wire g5477A;
wire g6910A;
wire g10417A;
wire I15986A;
wire g713A;
wire g2237A;
wire g6488A;
wire g7712A;
wire g7897A;
wire g6828A;
wire g7638A;
wire g3015A;
wire g3121A;
wire I4917A;
wire g10800A;
wire g4300A;
wire g5420A;
wire g8019A;
wire I15956A;
wire g1840A;
wire g2557A;
wire g105A;
wire g9097A;
wire g6821A;
wire g3938A;
wire I5245A;
wire g253A;
wire g7682A;
wire g8267A;
wire g11478A;
wire g3698A;
wire g4379A;
wire g4144A;
wire g584A;
wire g131A;
wire g2254A;
wire g4289A;
wire g3992A;
wire g4777A;
wire I5424A;
wire g1776A;
wire g4585A;
wire g7934A;
wire g8089A;
wire g243A;
wire g2438A;
wire g6516A;
wire g8244A;
wire g4271A;
wire g4753A;
wire g8631A;
wire g4807A;
wire g10793A;
wire g7045A;
wire g5910A;
wire g9454A;
wire g686A;
wire g2212A;
wire I14299A;
wire g2563A;
wire g3141A;
wire g2478A;
wire g569A;
wire g35A;
wire g3215A;
wire g3710A;
wire I16252A;
wire g10726A;
wire g7516A;
wire g7920A;
wire g6824A;
wire g162A;
wire g2229A;
wire g9931A;
wire I15157A;
wire g11157A;
wire I15365A;
wire g79A;
wire I9279A;
wire g5361A;
wire g10558A;
wire g5248A;
wire g3880A;
wire g5557A;
wire g2172A;
wire g6759A;
wire g6502A;
wire g10797A;
wire g8241A;
wire I5044A;
wire g7685A;
wire g4471A;
wire g10780A;
wire g11625A;
wire g11372A;
wire g10007A;
wire I15287A;
wire g10771A;
wire I15290A;
wire g9720A;
wire g127A;
wire g2249A;
wire g5803A;
wire g11231A;
wire g11580A;
wire g5478A;
wire g11243A;
wire g4998A;
wire g10019A;
wire I5414A;
wire g4114A;
wire g11293A;
wire g2176A;
wire g4779A;
wire g5820A;
wire g8173A;
wire g3111A;
wire g3628A;
wire g4977A;
wire g6081A;
wire g255A;
wire g6533A;
wire I8503A;
wire g7460A;
wire g7910A;
wire g1984A;
wire g3688A;
wire g4285A;
wire g5867A;
wire g6354A;
wire g1690A;
wire g2031A;
wire g1857A;
wire I5510A;
wire g10405A;
wire g7932A;
wire g8085A;
wire g928A;
wire g7883A;
wire g10448A;
wire g5001A;
wire g8245A;
wire g3440A;
wire g4737A;
wire g8451A;
wire g8214A;
wire I13351A;
wire g3041A;
wire g10767A;
wire g10599A;
wire g10501A;
wire g3546A;
wire g8512A;
wire g2276A;
wire g6000A;
wire g6863A;
wire g10809A;
wire g10883A;
wire g5521A;
wire I14323A;
wire g11492A;
wire g932A;
wire g37A;
wire I6260A;
wire I9311A;
wire g4490A;
wire g8488A;
wire I5579A;
wire I9268A;
wire g4903A;
wire g10720A;
wire g10334A;
wire g10439A;
wire g6934A;
wire g5309A;
wire g5878A;
wire g4273A;
wire g7622A;
wire g6123A;
wire g7467A;
wire g774A;
wire g1990A;
wire g2248A;
wire g6838A;
wire g2045A;
wire g4905A;
wire g10798A;
wire g10785A;
wire g8187A;
wire I13436A;
wire g605A;
wire g2399A;
wire g7204A;
wire g6830A;
wire g6716A;
wire g8944A;
wire I5254A;
wire g5543A;
wire I5410A;
wire g5300A;
wire g8921A;
wire g8745A;
wire g8849A;
wire g6096A;
wire I7752A;
wire g6003A;
wire g3431A;
wire I7840A;
wire g10852A;
wire g6733A;
wire g7562A;
wire g6548A;
wire g1419A;
wire I9810A;
wire g5502A;
wire g260A;
wire g4679A;
wire g6823A;
wire g4890A;
wire g7981A;
wire g2579A;
wire g3776A;
wire g572A;
wire g3381A;
wire g10863A;
wire g971A;
wire g2008A;
wire g8039A;
wire g6526A;
wire g1900A;
wire g2336A;
wire g10664A;
wire g7189A;
wire g5278A;
wire g8923A;
wire g5173A;
wire g3521A;
wire I14306A;
wire g10712A;
wire I9296A;
wire g4264A;
wire g2178A;
wire g6755A;
wire g2791A;
wire I6962A;
wire g5226A;
wire g704A;
wire g2230A;
wire g4437A;
wire g11514A;
wire g7505A;
wire g38A;
wire g9507A;
wire g10411A;
wire I15974A;
wire g4506A;
wire g1834A;
wire g2550A;
wire g10348A;
wire g10400A;
wire I9282A;
wire I5584A;
wire g9324A;
wire g3664A;
wire g10001A;
wire g5526A;
wire g7697A;
wire g231A;
wire g2395A;
wire I5395A;
wire g4788A;
wire g4465A;
wire g8289A;
wire g6403A;
wire g8203A;
wire I15510A;
wire g5403A;
wire g6902A;
wire g6015A;
wire g11340A;
wire g6542A;
wire I5406A;
wire g3744A;
wire g581A;
wire I4883A;
wire g4537A;
wire g7688A;
wire g882A;
wire g2481A;
wire g6507A;
wire g10485A;
wire I4935A;
wire g10683A;
wire I9308A;
wire I5070A;
wire g5556A;
wire g8505A;
wire g8603A;
wire g11641A;
wire g3423A;
wire g4787A;
wire I9332A;
wire g10765A;
wire g6447A;
wire g4801A;
wire g11305A;
wire g3092A;
wire g6126A;
wire g4281A;
wire g5493A;
wire g5613A;
wire g639A;
wire g10414A;
wire g7986A;
wire g8255A;
wire g8000A;
wire g8081A;
wire g814A;
wire I9479A;
wire I4780A;
wire g2216A;
wire g10522A;
wire I5383A;
wire g8060A;
wire g7191A;
wire g8746A;
wire g8783A;
wire g10557A;
wire g5150A;
wire I5445A;
wire g4449A;
wire I4866A;
wire g6469A;
wire g7696A;
wire g10452A;
wire g4498A;
wire g8744A;
wire g8828A;
wire g2034A;
wire g2677A;
wire g5514A;
wire g6627A;
wire g4893A;
wire g10268A;
wire g10361A;
wire g3737A;
wire g9257A;
wire g9525A;
wire g5194A;
wire g668A;
wire g2198A;
wire g3418A;
wire I7771A;
wire g6901A;
wire g8043A;
wire g5263A;
wire g6929A;
wire g5857A;
wire g3523A;
wire g8049A;
wire g4529A;
wire g9699A;
wire g722A;
wire g2241A;
wire g6786A;
wire g7218A;
wire g7681A;
wire g6234A;
wire g5824A;
wire g7101A;
wire g10864A;
wire g7651A;
wire g7914A;
wire g986A;
wire I13427A;
wire g8816A;
wire I14319A;
wire I5430A;
wire g2175A;
wire g10862A;
wire I15980A;
wire g11077A;
wire I9259A;
wire g7683A;
wire I16717A;
wire I5388A;
wire I9326A;
wire g153A;
wire g2211A;
wire g3222A;
wire g3983A;
wire g4678A;
wire g3101A;
wire g3543A;
wire I5053A;
wire g9268A;
wire g5942A;
wire g10331A;
wire g10421A;
wire g10721A;
wire g8051A;
wire g2118A;
wire g10383A;
wire g6541A;
wire g936A;
wire g9088A;
wire g139A;
wire g2083A;
wire I6360A;
wire g10773A;
wire g8193A;
wire I4992A;
wire g6523A;
wire I16982A;
wire g8546A;
wire g8599A;
wire g794A;
wire g1828A;
wire g2061A;
wire g746A;
wire g2187A;
wire I9383A;
wire g5404A;
wire g11393A;
wire g5258A;
wire g1845A;
wire g2271A;
wire g1400A;
wire g2446A;
wire g8265A;
wire g2984A;
wire g11561A;
wire g11575A;
wire g822A;
wire g4765A;
wire g4334A;
wire g1936A;
wire g2345A;
wire g11233A;
wire g7950A;
wire g8106A;
wire g6586A;
wire g6908A;
wire g8768A;
wire g8885A;
wire g563A;
wire g33A;
wire g5808A;
wire I5418A;
wire g1361A;
wire g2016A;
wire g5271A;
wire g6333A;
wire g10515A;
wire g7692A;
wire I9273A;
wire g6045A;
wire g123A;
wire g731A;
wire g2251A;
wire g1988A;
wire g2047A;
wire g10927A;
wire g7590A;
wire g2275A;
wire g6468A;
wire g10782A;
wire g10886A;
wire g6672A;
wire g6840A;
wire g5230A;
wire g549A;
wire g8743A;
wire g8858A;
wire g3354A;
wire g4671A;
wire g5914A;
wire g7705A;
wire g7953A;
wire g8115A;
wire g10025A;
wire g1218A;
wire g2017A;
wire I5101A;
wire g6038A;
wire g1882A;
wire g2328A;
wire I5057A;
wire g1868A;
wire g2542A;
wire g4488A;
wire g1891A;
wire g2330A;
wire g3863A;
wire g6471A;
wire g11303A;
wire I9276A;
wire g7949A;
wire I5041A;
wire g782A;
wire g1992A;
wire I5441A;
wire g1110A;
wire g4365A;
wire g5266A;
wire g8234A;
wire I13364A;
wire g4158A;
wire g10663A;
wire g8920A;
wire g4283A;
wire I4859A;
wire g10788A;
wire g1397A;
wire g2456A;
wire g7512A;
wire g7919A;
wire g4484A;
wire I17413A;
wire I9346A;
wire g643A;
wire g1976A;
wire g7952A;
wire g865A;
wire I4820A;
wire I5435A;
wire g8815A;
wire I14315A;
wire g3008A;
wire g4467A;
wire g9713A;
wire g4290A;
wire g7527A;
wire g4770A;
wire g9474A;
wire g36A;
wire g5842A;
wire I9265A;
wire g7671A;
wire g8056A;
wire g8700A;
wire g4381A;
wire g5396A;
wire g1854A;
wire g7203A;
wire I6273A;
wire g10382A;
wire g10583A;
wire g10629A;
wire g8045A;
wire g7843A;
wire g2652A;
wire g754A;
wire g2057A;
wire g3539A;
wire g4263A;
wire g8269A;
wire I9349A;
wire I13323A;
wire g1386A;
wire g2549A;
wire g5261A;
wire g3104A;
wire g3419A;
wire g3425A;
wire I7829A;
wire g9802A;
wire g806A;
wire g6537A;
wire I13338A;
wire g5221A;
wire g3086A;
wire g2253A;
wire g4902A;
wire g6080A;
wire I9371A;
wire g5485A;
wire g6059A;
wire g4089A;
wire I5588A;
wire g7664A;
wire g7907A;
wire g4673A;
wire g8551A;
wire g5126A;
wire g10866A;
wire g10597A;
wire g11603A;
wire g6332A;
wire g4231A;
wire g9526A;
wire g207A;
wire g2570A;
wire g7473A;
wire g7915A;
wire I4783A;
wire g1991A;
wire g7677A;
wire g64A;
wire g11249A;
wire g636A;
wire g2506A;
wire g11348A;
wire g10779A;
wire g11488A;
wire g3491A;
wire g40A;
wire g3438A;
wire I7852A;
wire g757A;
wire g5354A;
wire g5295A;
wire g5918A;
wire g6894A;
wire g3513A;
wire g1713A;
wire I6240A;
wire g258A;
wire g591A;
wire g2374A;
wire g9424A;
wire g4076A;
wire g6534A;
wire g58A;
wire g3793A;
wire g6928A;
wire g7686A;
wire g3414A;
wire I7825A;
wire g8055A;
wire g11291A;
wire g237A;
wire g2420A;
wire g3209A;
wire g4739A;
wire g5509A;
wire g6833A;
wire g1958A;
wire g6918A;
wire g4608A;
wire I4948A;
wire g6915A;
wire g6911A;
wire I5060A;
wire g8812A;
wire I9237A;
wire g4553A;
wire g7441A;
wire g5996A;
wire g8047A;
wire g1786A;
wire g6653A;
wire g7438A;
wire g6832A;
wire I5047A;
wire g4771A;
wire g11481A;
wire g10857A;
wire g7947A;
wire g8100A;
wire g3681A;
wire g7918A;
wire I5427A;
wire g6478A;
wire g4117A;
wire g6897A;
wire g6042A;
wire I9717A;
wire g119A;
wire g11229A;
wire g1453A;
wire g2410A;
wire g10402A;
wire g4342A;
wire g4330A;
wire g8221A;
wire g1927A;
wire g2343A;
wire g11609A;
wire g10859A;
wire g6054A;
wire g6508A;
wire g6531A;
wire g8050A;
wire g8261A;
wire I9290A;
wire g11376A;
wire g580A;
wire I4876A;
wire g802A;
wire g8559A;
wire I9769A;
wire g2260A;
wire g10556A;
wire g148A;
wire g2202A;
wire g7032A;
wire g8390A;
wire g8548A;
wire g590A;
wire g2518A;
wire g4548A;
wire g4293A;
wire I16507A;
wire g5390A;
wire g4561A;
wire g8233A;
wire g1289A;
wire g8200A;
wire g4294A;
wire g76A;
wire g8767A;
wire g3071A;
wire g3723A;
wire I15962A;
wire g940A;
wire g7987A;
wire g8094A;
wire g1861A;
wire g2050A;
wire g1987A;
wire g4480A;
wire g11483A;
wire g1351A;
wire g10702A;
wire g5863A;
wire g2273A;
wire g5392A;
wire g9082A;
wire g5838A;
wire g8270A;
wire g10776A;
wire g2024A;
wire g2777A;
wire g6513A;
wire g9272A;
wire g10732A;
wire g1411A;
wire g10898A;
wire g869A;
wire g8052A;
wire g4325A;
wire g3368A;
wire g762A;
wire g4421A;
wire I8869A;
wire g5319A;
wire g8766A;
wire g10555A;
wire g586A;
wire g61A;
wire g6205A;
wire g778A;
wire g622A;
wire g8820A;
wire I9329A;
wire g11199A;
wire g9124A;
wire g6839A;
wire g6522A;
wire g10936A;
wire g7852A;
wire g7923A;
wire g11320A;
wire g6841A;
wire g10328A;
wire g10431A;
wire g8769A;
wire g6224A;
wire g2208A;
wire g11349A;
wire g4782A;
wire g6470A;
wire g11225A;
wire g5755A;
wire g4292A;
wire g1212A;
wire g6515A;
wire g3003A;
wire g3760A;
wire g9710A;
wire g5117A;
wire g3631A;
wire g5182A;
wire g11430A;
wire I9368A;
wire g10791A;
wire g5004A;
wire g1806A;
wire g7632A;
wire g11485A;
wire I5399A;
wire g6331A;
wire g1718A;
wire g2424A;
wire g5257A;
wire g8053A;
wire g4518A;
wire g7550A;
wire g219A;
wire g2077A;
wire g3103A;
wire g4764A;
wire g7913A;
wire g1989A;
wire g3068A;
wire g6109A;
wire I15500A;
wire g5763A;
wire g6480A;
wire g6795A;
wire g6449A;
wire g8194A;
wire g2257A;
wire g5201A;
wire g5269A;
wire g7497A;
wire g876A;
wire g2444A;
wire g1107A;
wire g8938A;
wire g7990A;
wire g8099A;
wire g4238A;
wire g8775A;
wire g4891A;
wire g8266A;
wire g11290A;
wire g6501A;
wire g10570A;
wire g10676A;
wire g6334A;
wire g786A;
wire g1993A;
wire g10719A;
wire g1104A;
wire g4727A;
wire g4274A;
wire g8765A;
wire g6916A;
wire g8811A;
wire I14303A;
wire g5174A;
wire I5525A;
wire I14330A;
wire g583A;
wire I4900A;
wire g11308A;
wire g3060A;
wire g5847A;
wire g10554A;
wire g10784A;
wire g2979A;
wire g599A;
wire g2382A;
wire g7680A;
wire g10396A;
wire g3784A;
wire g11425A;
wire I14295A;
wire g1346A;
wire I9293A;
wire I5815A;
wire g4002A;
wire g7062A;
wire g3479A;
wire g5548A;
wire g6131A;
wire g2449A;
wire g6820A;
wire g3390A;
wire g5627A;
wire g3501A;
wire g4340A;
wire I13385A;
wire g143A;
wire g2095A;
wire g1771A;
wire g257A;
wire g2297A;
wire g262A;
wire g6922A;
wire g1969A;
wire g6747A;
wire g11391A;
wire g8818A;
wire g8649A;
wire g9555A;
wire g6071A;
wire g1796A;
wire g7942A;
wire g8095A;
wire g6718A;
wire g611A;
wire g2364A;
wire g10858A;
wire g55A;
wire g1864A;
wire g2054A;
wire g2018A;
wire g2725A;
wire g627A;
wire g8926A;
wire g4239A;
wire g11602A;
wire g8041A;
wire g5503A;
wire g646A;
wire g1980A;
wire g981A;
wire g8164A;
wire g883A;
wire I6220A;
wire g582A;
wire I4891A;
wire g8922A;
wire g5536A;
wire g578A;
wire g5810A;
wire g7067A;
wire g8236A;
wire g11605A;
wire g8048A;
wire g6528A;
wire g1909A;
wire g2338A;
wire g34A;
wire g6524A;
wire g7446A;
wire g3056A;
wire g3475A;
wire g7258A;
wire g7219A;
wire g8046A;
wire g3706A;
wire g4822A;
wire g11482A;
wire g10381A;
wire g4477A;
wire g10333A;
wire g10437A;
wire g4456A;
wire g2310A;
wire g3039A;
wire g6923A;
wire g4255A;
wire g878A;
wire g790A;
wire g4732A;
wire g8937A;
wire g4752A;
wire g6538A;
wire g10339A;
wire g3524A;
wire g11306A;
wire g7183A;
wire g4778A;
wire g6165A;
wire g6895A;
wire g588A;
wire g11223A;
wire g6163A;
wire g6179A;
wire g9052A;
wire g9505A;
wire g9721A;
wire g654A;
wire g2268A;
wire g8776A;
wire g6827A;
wire g461A;
wire g4309A;
wire g9331A;
wire g7244A;
wire g7586A;
wire g7930A;
wire g5222A;
wire g11300A;
wire g10718A;
wire g213A;
wire g2070A;
wire g3906A;
wire g579A;
wire g5445A;
wire g11227A;
wire g6088A;
wire g658A;
wire g2331A;
wire g1365A;
wire g2406A;
wire g8206A;
wire I13332A;
wire g6679A;
wire g11636A;
wire g11239A;
wire g11219A;
wire g225A;
wire g2087A;
wire g2117A;
wire g2801A;
wire g3062A;
wire g3738A;
wire g9266A;
wire g9760A;
wire g11608A;
wire g8059A;
wire g8771A;
wire g2459A;
wire g6035A;
wire g1811A;
wire g7106A;
wire g471A;
wire g6198A;
wire g7992A;
wire g8105A;
wire g2169A;
wire g8973A;
wire g617A;
wire g2369A;
wire g6834A;
wire g197A;
wire g2407A;
wire g1962A;
wire g5148A;
wire I14642A;
wire g5836A;
wire g7134A;
wire I15514A;
wire g10795A;
wire g11083A;
wire g11276A;
wire g10770A;
wire g1810A;
wire g9271A;
wire g677A;
wire g2203A;
wire g587A;
wire I5497A;
wire I13421A;
wire g10494A;
wire g8773A;
wire g3462A;
wire I16220A;
wire g3662A;
wire g6740A;
wire g10484A;
wire g7143A;
wire g8939A;
wire g1703A;
wire g2028A;
wire g8772A;
wire g4336A;
wire g2067A;
wire g1814A;
wire g2564A;
wire g6093A;
wire g6500A;
wire g1407A;
wire g3705A;
wire g10500A;
wire g2794A;
wire g4065A;
wire g4243A;
wire g4934A;
wire g6485A;
wire g8777A;
wire g6244A;
wire g5304A;
wire g11640A;
wire g3814A;
wire g4784A;
wire g11487A;
wire g9110A;
wire g1822A;
wire g2571A;
wire g11380A;
wire g1950A;
wire g826A;
wire g9269A;
wire g7054A;
wire g1975A;
wire g7236A;
wire g2774A;
wire g3247A;
wire g3967A;
wire g11314A;
wire g585A;
wire g5276A;
wire g9150A;
wire g1389A;
wire g2396A;
wire g11298A;
wire g7202A;
wire g6819A;
wire g2987A;
wire g758A;
wire g11539A;
wire g1336A;
wire g108A;
wire g5317A;
wire g67A;
wire g10453A;
wire g6243A;
wire g6514A;
wire g8817A;
wire g8810A;
wire g1206A;
wire I6277A;
wire g1368A;
wire g2381A;
wire g9313A;
wire g10387A;
wire g6983A;
wire g8366A;
wire g8509A;
wire g7450A;
wire g7905A;
wire g4473A;
wire g6577A;
wire g1341A;
wire g1374A;
wire g2421A;
wire g3200A;
wire g4001A;
wire g8040A;
wire g5255A;
wire g6900A;
wire g8042A;
wire g11490A;
wire g11515A;
wire g8230A;
wire g6546A;
wire g3485A;
wire g1383A;
wire g2562A;
wire g6697A;
wire g8574A;
wire g5770A;
wire I11360A;
wire g8889A;
wire g10711A;
wire g9719A;
wire g11312A;
wire g5287A;
wire g11107A;
wire g1791A;
wire g6351A;
wire g9778A;
wire g6479A;
wire g3120A;
wire g3765A;
wire g5814A;
wire g5849A;
wire g1101A;
wire g575A;
wire g10559A;
wire g5219A;
wire g7240A;
wire I9352A;
wire g8819A;
wire g9256A;
wire g261A;
wire g6656A;
wire g976A;
wire g736A;
wire g1424A;
wire g1377A;
wire g2074A;
wire g6906A;
wire g10717A;
wire g4759A;
wire g5189A;
wire g8770A;
wire g6392A;
wire g6621A;
wire g11610A;
wire g4582A;
wire g6432A;
wire g7454A;
wire g7908A;
wire g8264A;
wire g11604A;
wire g9764A;
wire g2161A;
wire g3291A;
wire g7245A;
wire g2510A;
wire g256A;
wire g2439A;
wire g3207A;
wire g810A;
wire g11486A;
wire g12A;
wire g2126A;
wire g7581A;
wire g10799A;
wire I15507A;
wire I9221A;
wire g114A;
wire g1964A;
wire g10357A;
wire g6439A;
wire g8507A;
wire g8688A;
wire g7133A;
wire g8642A;
wire g8044A;
wire g8254A;
wire g11549A;
wire g1357A;
wire g2023A;
wire g7379A;
wire g11232A;
wire g11607A;
wire g6573A;
wire g3506A;
wire g3407A;
wire g770A;
wire g6193A;
wire g3108A;
wire g3408A;
wire g248A;
wire g2451A;
wire g7225A;
wire g8220A;
wire g7231A;
wire g4576A;
wire g3943A;
wire g4904A;
wire g8806A;
wire g11292A;
wire g6822A;
wire g7624A;
wire g3661A;
wire I15861A;
wire g73A;
wire g1801A;
wire g8327A;
wire g6912A;
wire g6898A;
wire g554A;
wire g8146A;
wire I5020A;
wire g5421A;
wire g1766A;
wire g7994A;
wire g8103A;
wire g1362A;
wire g2434A;
wire g3913A;
wire g6702A;
wire g4880A;
wire g8696A;
wire g868A;
wire g8813A;
wire I14309A;
wire g1945A;
wire g2347A;
wire g6924A;
wire g5308A;
wire g7574A;
wire g11310A;
wire g11294A;
wire g5852A;
wire g2970A;
wire g6026A;
wire g10369A;
wire g5286A;
wire g4554A;
wire g8024A;
wire g8945A;
wire g4804A;
wire g6525A;
wire g1380A;
wire g2060A;
wire g6019A;
wire g6617A;
wire g8210A;
wire g5083A;
wire g3585A;
wire g589A;
wire g7541A;
wire g4760A;
wire g26A;
wire g2479A;
wire g10860A;
wire g10502A;
wire g11579A;
wire g11639A;
wire g9814A;
wire g5030A;
wire g39A;
wire g6826A;
wire g2303A;
wire g9773A;
wire g52A;
wire g7626A;
wire g5200A;
wire g4457A;
wire g6829A;
wire g7211A;
wire g466A;
wire g456A;
wire g7660A;
wire g10722A;
wire g8887A;
wire g11484A;
wire g11286A;
wire g6002A;
wire g11606A;
wire g11217A;
wire g10454A;
wire g6757A;
wire g6216A;
wire g8941A;
wire g10856A;
wire g4892A;
wire g7903A;
wire g6930A;
wire g8250A;
wire g5250A;
wire g4525A;
wire g6049A;
wire g8943A;
wire g10861A;
wire g192A;
wire g2475A;
wire g8779A;
wire g766A;
wire g5484A;
wire g557A;
wire g11203A;
wire g3304A;
wire g6557A;
wire g4482A;
wire g1781A;
wire g5190A;
wire g6180A;
wire g5274A;
wire g8774A;
wire g10325A;
wire g10444A;
wire g566A;
wire g8260A;
wire g6099A;
wire g10401A;
wire g6831A;
wire g6068A;
wire g7137A;
wire g7917A;
wire g9473A;
wire g1965A;
wire g6545A;
wire g11547A;
wire g7257A;
wire g6909A;
wire g8384A;
wire g1872A;
wire g2503A;
wire g11392A;
wire g6506A;
wire g8883A;
wire g695A;
wire g2224A;
wire g6728A;
wire g10724A;
wire g4556A;
wire g3070A;
wire g2250A;
wire g11103A;
wire g9900A;
wire g845A;
wire g11095A;
wire g1645A;
wire g4973A;
wire g7389A;
wire g7465A;
wire g7888A;
wire g1642A;
wire g4969A;
wire g8224A;
wire g2892A;
wire g5686A;
wire g10308A;
wire g4123A;
wire g8120A;
wire g287A;
wire g6788A;
wire g4824A;
wire g5598A;
wire g278A;
wire g9694A;
wire g10495A;
wire g1684A;
wire g2945A;
wire g11190A;
wire g8639A;
wire g8789A;
wire g9728A;
wire g9563A;
wire g9852A;
wire g1053A;
wire g5625A;
wire g995A;
wire g4875A;
wire g1574A;
wire g9701A;
wire g7138A;
wire g10752A;
wire g11058A;
wire g11211A;
wire g435A;
wire g11024A;
wire g8307A;
wire g8547A;
wire g10669A;
wire g691A;
wire g7707A;
wire g3813A;
wire g4884A;
wire g4839A;
wire g1561A;
wire g9870A;
wire g6640A;
wire g9240A;
wire g9650A;
wire g5687A;
wire g7957A;
wire g3512A;
wire g7449A;
wire g1011A;
wire g4235A;
wire g345A;
wire g4343A;
wire g11296A;
wire g1A;
wire g9292A;
wire g9594A;
wire g1160A;
wire g9923A;
wire g9367A;
wire g9943A;
wire g1721A;
wire g5525A;
wire g440A;
wire g8876A;
wire g476A;
wire g10564A;
wire g10705A;
wire g9913A;
wire g9624A;
wire g9934A;
wire g6225A;
wire g1240A;
wire g6324A;
wire g10686A;
wire g1223A;
wire g6540A;
wire g8663A;
wire g1308A;
wire g11581A;
wire g6206A;
wire g452A;
wire g3989A;
wire g7260A;
wire g7730A;
wire g1235A;
wire g7504A;
wire g1887A;
wire g7185A;
wire I5689A;
wire I5690A;
wire g7881A;
wire g11070A;
wire g9736A;
wire g9859A;
wire g8877A;
wire g2274A;
wire g11590A;
wire g6199A;
wire g8932A;
wire g1730A;
wire g5545A;
wire g5180A;
wire g1615A;
wire g5591A;
wire g8412A;
wire g8556A;
wire g374A;
wire g11094A;
wire g5044A;
wire g5853A;
wire g6245A;
wire g4360A;
wire g8930A;
wire g5507A;
wire g3087A;
wire g11150A;
wire g8302A;
wire g8464A;
wire g272A;
wire g9692A;
wire g1428A;
wire g4996A;
wire g7131A;
wire g421A;
wire g11019A;
wire g9951A;
wire g9536A;
wire g9960A;
wire g11196A;
wire g11018A;
wire g10550A;
wire g10595A;
wire g10433A;
wire g10544A;
wire g10623A;
wire g4878A;
wire g4838A;
wire g5204A;
wire g8609A;
wire g8844A;
wire g6185A;
wire g6701A;
wire g10725A;
wire g5100A;
wire g1089A;
wire g4882A;
wire g8731A;
wire g1504A;
wire g5128A;
wire g1932A;
wire g6886A;
wire g8415A;
wire g8557A;
wire g8966A;
wire g8071A;
wire g11597A;
wire g9722A;
wire g9785A;
wire g9828A;
wire g1672A;
wire g2918A;
wire g9725A;
wire g9830A;
wire g8955A;
wire g4A;
wire g9592A;
wire g1618A;
wire g5123A;
wire g6078A;
wire g7059A;
wire g7459A;
wire g861A;
wire g11102A;
wire g709A;
wire g7718A;
wire g7535A;
wire g1577A;
wire g9703A;
wire g5528A;
wire g9911A;
wire g9932A;
wire g1636A;
wire g5530A;
wire g2760A;
wire g8629A;
wire g6187A;
wire g6887A;
wire g5605A;
wire g6228A;
wire g1275A;
wire g6322A;
wire I6337A;
wire I6338A;
wire g8967A;
wire g1458A;
wire g5010A;
wire g3275A;
wire g1678A;
wire g2895A;
wire g7721A;
wire g1549A;
wire g9866A;
wire g1534A;
wire g9716A;
wire g10744A;
wire g10808A;
wire g1231A;
wire g3047A;
wire g3685A;
wire g4492A;
wire g8614A;
wire g8822A;
wire g10560A;
wire g11456A;
wire g9724A;
wire g9848A;
wire g4714A;
wire g6550A;
wire g5172A;
wire g10642A;
wire g2531A;
wire g3284A;
wire g284A;
wire g302A;
wire g9855A;
wire g1630A;
wire g5618A;
wire g6891A;
wire g7940A;
wire g312A;
wire g11085A;
wire g396A;
wire g1432A;
wire g4968A;
wire g8646A;
wire g8837A;
wire g9125A;
wire g9644A;
wire g1546A;
wire g5804A;
wire g8300A;
wire g8462A;
wire I6330A;
wire g333A;
wire g11156A;
wire g293A;
wire g6342A;
wire g1552A;
wire g9867A;
wire g1537A;
wire g9717A;
wire g4871A;
wire g10435A;
wire g426A;
wire g7741A;
wire g1327A;
wire g9151A;
wire g9386A;
wire g8607A;
wire g8842A;
wire g8A;
wire g9599A;
wire g8974A;
wire g9274A;
wire g5518A;
wire g9111A;
wire g9614A;
wire g4122A;
wire g4610A;
wire g7217A;
wire g11557A;
wire g1675A;
wire g2911A;
wire g11210A;
wire g7466A;
wire g9918A;
wire g9939A;
wire g11279A;
wire g10513A;
wire g10440A;
wire I16145A;
wire g10518A;
wire g1129A;
wire g7055A;
wire g1095A;
wire g5264A;
wire g1265A;
wire g6329A;
wire g8176A;
wire g7510A;
wire g8005A;
wire g3281A;
wire g4099A;
wire g11601A;
wire g11187A;
wire g6746A;
wire g6221A;
wire g8630A;
wire g9622A;
wire g10923A;
wire g11143A;
wire g9886A;
wire g9676A;
wire g9904A;
wire g8733A;
wire g348A;
wire g6624A;
wire g530A;
wire g11169A;
wire g8073A;
wire g9706A;
wire g9512A;
wire g9841A;
wire g5592A;
wire g5882A;
wire g8645A;
wire g8796A;
wire g534A;
wire g11168A;
wire g1015A;
wire g4269A;
wire g727A;
wire g1047A;
wire g5611A;
wire g673A;
wire g8069A;
wire g1567A;
wire g9695A;
wire g10304A;
wire g8305A;
wire g8469A;
wire g1071A;
wire g4712A;
wire g5762A;
wire g6576A;
wire g10622A;
wire g5217A;
wire g11015A;
wire g5674A;
wire g9173A;
wire g9359A;
wire g8960A;
wire g9223A;
wire g11556A;
wire g1595A;
wire g9858A;
wire g5541A;
wire g363A;
wire g4534A;
wire g1499A;
wire g5897A;
wire g6177A;
wire g6699A;
wire g6855A;
wire g3098A;
wire g3804A;
wire g5680A;
wire g9642A;
wire g1528A;
wire g5744A;
wire g8399A;
wire g1762A;
wire g9030A;
wire g9447A;
wire g1849A;
wire g516A;
wire g11178A;
wire g8414A;
wire g8510A;
wire g1296A;
wire g6319A;
wire g11186A;
wire g1681A;
wire g2951A;
wire g6352A;
wire g9205A;
wire g9595A;
wire g4109A;
wire g4831A;
wire g1654A;
wire g5492A;
wire g8934A;
wire g10312A;
wire g6186A;
wire g9612A;
wire g1738A;
wire g9417A;
wire g9914A;
wire g9935A;
wire g10658A;
wire g10745A;
wire g956A;
wire g11216A;
wire g8971A;
wire g9328A;
wire g11587A;
wire g1245A;
wire g6325A;
wire g431A;
wire g7368A;
wire g552A;
wire g6083A;
wire g1227A;
wire g6544A;
wire g5476A;
wire g7743A;
wire g1083A;
wire g4869A;
wire g1598A;
wire g5722A;
wire g5813A;
wire g6790A;
wire g8408A;
wire g10761A;
wire g7734A;
wire g7926A;
wire g8136A;
wire g5569A;
wire g401A;
wire g9392A;
wire g9902A;
wire g8623A;
wire g1657A;
wire g5500A;
wire g2496A;
wire g3010A;
wire g5877A;
wire g6756A;
wire g8972A;
wire g336A;
wire g6622A;
wire g11612A;
wire g1311A;
wire g9366A;
wire g11230A;
wire g1284A;
wire g1215A;
wire g4364A;
wire g9649A;
wire g1543A;
wire g5795A;
wire g1524A;
wire g5737A;
wire g1753A;
wire g4054A;
wire g5823A;
wire g6345A;
wire g11275A;
wire g296A;
wire g9851A;
wire g5802A;
wire g6763A;
wire g416A;
wire g10511A;
wire g10509A;
wire g10507A;
wire I16142A;
wire g1571A;
wire g9698A;
wire g1032A;
wire g4725A;
wire g9954A;
wire g9964A;
wire g1663A;
wire g5523A;
wire g8402A;
wire g8550A;
wire g8611A;
wire g8845A;
wire g2081A;
wire g281A;
wire g6359A;
wire g1324A;
wire g11586A;
wire g5147A;
wire g11007A;
wire g5104A;
wire g4821A;
wire g5099A;
wire g5919A;
wire g1627A;
wire g5499A;
wire g3529A;
wire g4389A;
wire g3497A;
wire g6416A;
wire g1444A;
wire g4990A;
wire g9010A;
wire g9619A;
wire I6630A;
wire g6047A;
wire g953A;
wire g9652A;
wire g10505A;
wire g10469A;
wire g9711A;
wire g9519A;
wire g9843A;
wire g1074A;
wire g5273A;
wire g11465A;
wire g4348A;
wire g11237A;
wire g9731A;
wire g9834A;
wire g6654A;
wire g1041A;
wire g5444A;
wire g3714A;
wire g11285A;
wire g9598A;
wire g8097A;
wire g8726A;
wire g4816A;
wire g6880A;
wire g1157A;
wire g3287A;
wire g10759A;
wire g9917A;
wire g9938A;
wire g10652A;
wire g10758A;
wire g406A;
wire g9891A;
wire g9909A;
wire g6663A;
wire g7127A;
wire g11165A;
wire g1260A;
wire g6328A;
wire g8401A;
wire g5125A;
wire g11006A;
wire g1080A;
wire g4865A;
wire g1077A;
wire g4715A;
wire g2325A;
wire g4604A;
wire g5513A;
wire g965A;
wire g11222A;
wire g1145A;
wire g6554A;
wire g7732A;
wire g9586A;
wire g4401A;
wire g4104A;
wire g5178A;
wire g4584A;
wire g7472A;
wire g11253A;
wire g9860A;
wire g11600A;
wire g1586A;
wire g9645A;
wire g11236A;
wire g3106A;
wire g4162A;
wire g553A;
wire g6090A;
wire g269A;
wire g9691A;
wire g11316A;
wire g501A;
wire g11175A;
wire g664A;
wire g8068A;
wire g9607A;
wire g9952A;
wire g9962A;
wire g6348A;
wire g9659A;
wire g1318A;
wire g9358A;
wire I6316A;
wire I6317A;
wire g1711A;
wire g4486A;
wire g8995A;
wire g9587A;
wire g5632A;
wire g8965A;
wire g991A;
wire g4881A;
wire g11209A;
wire g8715A;
wire g8848A;
wire g3263A;
wire g4070A;
wire g6463A;
wire g1896A;
wire g7820A;
wire g448A;
wire g11021A;
wire g1044A;
wire g5917A;
wire g6619A;
wire g1300A;
wire g6318A;
wire g6872A;
wire g11201A;
wire g10489A;
wire g10514A;
wire g4006A;
wire g299A;
wire g9853A;
wire g11274A;
wire g8119A;
wire g1747A;
wire g9420A;
wire g5233A;
wire g7092A;
wire g6549A;
wire g11464A;
wire g4487A;
wire g1687A;
wire g2939A;
wire g6739A;
wire g7060A;
wire g1580A;
wire g5725A;
wire g11615A;
wire g2544A;
wire g11252A;
wire g5532A;
wire g3771A;
wire g11153A;
wire g9872A;
wire g9680A;
wire g9905A;
wire g7739A;
wire g6321A;
wire g8386A;
wire g8975A;
wire g2306A;
wire g6625A;
wire g7937A;
wire g8303A;
wire g8170A;
wire g5706A;
wire g2756A;
wire g8643A;
wire g8821A;
wire g5225A;
wire g10946A;
wire g4169A;
wire g5029A;
wire g11164A;
wire g4007A;
wire g1756A;
wire g4059A;
wire g1027A;
wire g4868A;
wire g5675A;
wire g4718A;
wire g10682A;
wire g6687A;
wire g682A;
wire g7704A;
wire g525A;
wire g1019A;
wire g4261A;
wire g3422A;
wire g5745A;
wire g8387A;
wire g7954A;
wire g11283A;
wire g8298A;
wire g8461A;
wire g10760A;
wire g11480A;
wire g6626A;
wire g6341A;
wire g10506A;
wire g16A;
wire g9648A;
wire g7453A;
wire g5995A;
wire g6645A;
wire g5707A;
wire g7548A;
wire g833A;
wire g11091A;
wire g496A;
wire g11174A;
wire g8403A;
wire g1250A;
wire g8605A;
wire g8841A;
wire g1914A;
wire g6879A;
wire g8763A;
wire g4502A;
wire g9702A;
wire g9839A;
wire g5841A;
wire g6358A;
wire g5575A;
wire g8107A;
wire g10240A;
wire g11192A;
wire g9618A;
wire g5539A;
wire g8416A;
wire g275A;
wire g9693A;
wire g11553A;
wire g7557A;
wire g1098A;
wire g5268A;
wire g9107A;
wire g10633A;
wire g7894A;
wire g8654A;
wire g9621A;
wire g5819A;
wire g6794A;
wire g3412A;
wire g7661A;
wire g2800A;
wire g3268A;
wire g9908A;
wire g3429A;
wire g351A;
wire g6628A;
wire g5470A;
wire g7526A;
wire g2204A;
wire g1482A;
wire g5025A;
wire g4921A;
wire g6204A;
wire g1750A;
wire g4048A;
wire g8935A;
wire g2525A;
wire g9593A;
wire g4827A;
wire g10701A;
wire g10733A;
wire g10777A;
wire g8130A;
wire g9955A;
wire g9965A;
wire g1710A;
wire g3684A;
wire g947A;
wire g11213A;
wire g1462A;
wire g5006A;
wire g9912A;
wire g9933A;
wire g8407A;
wire g8554A;
wire g9641A;
wire g6323A;
wire g10646A;
wire g10766A;
wire g6666A;
wire g4994A;
wire g5103A;
wire g3717A;
wire g11592A;
wire g1905A;
wire g6875A;
wire g9658A;
wire g6207A;
wire g6530A;
wire g8199A;
wire g7265A;
wire g9735A;
wire g9835A;
wire g6655A;
wire g3875A;
wire g7384A;
wire g7970A;
wire g1624A;
wire g5491A;
wire g8949A;
wire g11152A;
wire g9611A;
wire g2804A;
wire g6410A;
wire g10451A;
wire g4397A;
wire g5398A;
wire g7224A;
wire g5602A;
wire g6884A;
wire g8964A;
wire g11413A;
wire g1415A;
wire g4950A;
wire g5535A;
wire g6772A;
wire g7277A;
wire g8301A;
wire g8463A;
wire g2511A;
wire g10728A;
wire g6618A;
wire g6235A;
wire g6355A;
wire g3626A;
wire g4723A;
wire g8720A;
wire g6693A;
wire g11020A;
wire g1314A;
wire g11583A;
wire g8118A;
wire g8167A;
wire g7892A;
wire g8652A;
wire g5721A;
wire g10362A;
wire g10367A;
wire g9901A;
wire g290A;
wire g6792A;
wire g11282A;
wire g7945A;
wire g11302A;
wire g521A;
wire g3634A;
wire g11105A;
wire g8471A;
wire g8598A;
wire g7140A;
wire g9600A;
wire g1604A;
wire g9864A;
wire g11613A;
wire g5188A;
wire g7435A;
wire g7876A;
wire g1280A;
wire g4058A;
wire g5809A;
wire g6776A;
wire g630A;
wire g10301A;
wire g354A;
wire g4505A;
wire g17A;
wire g9623A;
wire g10739A;
wire g391A;
wire g11027A;
wire g10738A;
wire g8558A;
wire g8687A;
wire g6360A;
wire g1564A;
wire g9871A;
wire g5108A;
wire g11248A;
wire g4992A;
wire g11552A;
wire g944A;
wire g9651A;
wire g11204A;
wire g7824A;
wire g1133A;
wire g5115A;
wire g7102A;
wire g968A;
wire g9384A;
wire g2561A;
wire g9700A;
wire g9754A;
wire g9838A;
wire g10594A;
wire g10661A;
wire g11321A;
wire g8879A;
wire g7621A;
wire g8962A;
wire g2272A;
wire g10715A;
wire g8659A;
wire g950A;
wire g9643A;
wire g8957A;
wire g1669A;
wire g5538A;
wire g1744A;
wire g4000A;
wire g4126A;
wire g4088A;
wire g4400A;
wire I5886A;
wire I5887A;
wire g486A;
wire g6238A;
wire g10727A;
wire g8174A;
wire g305A;
wire g5067A;
wire g1512A;
wire g5418A;
wire g10297A;
wire g6353A;
wire g386A;
wire g11026A;
wire g11212A;
wire g4828A;
wire g6744A;
wire g1923A;
wire g10671A;
wire g2517A;
wire g4383A;
wire g4297A;
wire g5256A;
wire g4220A;
wire g8252A;
wire g8380A;
wire g7071A;
wire g9613A;
wire g8933A;
wire g5181A;
wire g7948A;
wire g324A;
wire g11149A;
wire g1601A;
wire g9862A;
wire g11387A;
wire g7955A;
wire g4161A;
wire g2321A;
wire g11148A;
wire g9712A;
wire g8931A;
wire g378A;
wire g11097A;
wire g3819A;
wire g2963A;
wire g11104A;
wire g1059A;
wire g6092A;
wire g4999A;
wire g4976A;
wire g632A;
wire g6858A;
wire g7409A;
wire g4103A;
wire I6309A;
wire g5944A;
wire g6580A;
wire g1056A;
wire g5631A;
wire g9414A;
wire g9660A;
wire g9926A;
wire g9946A;
wire I6331A;
wire g481A;
wire g9885A;
wire g9673A;
wire g9903A;
wire g10625A;
wire g6623A;
wire g11228A;
wire g11011A;
wire g1941A;
wire g6889A;
wire g7523A;
wire g7822A;
wire g8123A;
wire g11582A;
wire g4316A;
wire g3625A;
wire g10969A;
wire g5041A;
wire g9335A;
wire g9727A;
wire g9831A;
wire g9422A;
wire g4588A;
wire g8511A;
wire g8648A;
wire g8875A;
wire g5168A;
wire g7503A;
wire g7895A;
wire g8655A;
wire g1062A;
wire g4914A;
wire g9927A;
wire g9947A;
wire g1555A;
wire g5772A;
wire g1666A;
wire g5531A;
wire g5036A;
wire g10503A;
wire g7738A;
wire g8010A;
wire g8410A;
wire g5608A;
wire g6231A;
wire g10581A;
wire g10364A;
wire g10450A;
wire g2132A;
wire g2379A;
wire g9653A;
wire g1515A;
wire g10818A;
wire g8172A;
wire g10429A;
wire g5074A;
wire g1558A;
wire g9869A;
wire g10635A;
wire g10741A;
wire g8693A;
wire g5480A;
wire g3766A;
wire g4581A;
wire g2981A;
wire g8409A;
wire g8555A;
wire g9364A;
wire g506A;
wire g8994A;
wire g11299A;
wire g6592A;
wire g7958A;
wire g1474A;
wire g4995A;
wire g4079A;
wire g2264A;
wire g745A;
wire g2160A;
wire g3257A;
wire I6310A;
wire g1470A;
wire g5000A;
wire g3301A;
wire g1478A;
wire I5084A;
wire g1727A;
wire g9412A;
wire g1330A;
wire g9389A;
wire g10567A;
wire g10706A;
wire g10366A;
wire g10447A;
wire g10446A;
wire g10533A;
wire g5220A;
wire g10624A;
wire g10300A;
wire g5023A;
wire g4432A;
wire g4053A;
wire g7596A;
wire g1639A;
wire g5588A;
wire g6074A;
wire g9953A;
wire g9963A;
wire g3089A;
wire g3772A;
wire g5051A;
wire g8724A;
wire g4157A;
wire g1583A;
wire g9707A;
wire g8878A;
wire g10639A;
wire g10763A;
wire g6777A;
wire g8109A;
wire g7511A;
wire g7898A;
wire g11271A;
wire g11461A;
wire g5732A;
wire g315A;
wire g11145A;
wire g411A;
wire g11031A;
wire g1607A;
wire g9865A;
wire g1531A;
wire g9715A;
wire g9604A;
wire g8647A;
wire g8799A;
wire g11198A;
wire g6873A;
wire g6632A;
wire g6095A;
wire g9729A;
wire g9833A;
wire g1038A;
wire g6102A;
wire g7819A;
wire g11280A;
wire g7088A;
wire g9584A;
wire g9896A;
wire g8209A;
wire g6752A;
wire g11161A;
wire g8947A;
wire g5681A;
wire g7951A;
wire g9419A;
wire g1724A;
wire g5533A;
wire g8936A;
wire g178A;
wire g10670A;
wire g829A;
wire g11087A;
wire g4949A;
wire g5851A;
wire g6364A;
wire g7825A;
wire g1304A;
wire g10667A;
wire g7136A;
wire g339A;
wire g6532A;
wire g9385A;
wire g1436A;
wire g1440A;
wire g1448A;
wire g1137A;
wire g9897A;
wire g9425A;
wire g3383A;
wire g1035A;
wire g5601A;
wire g7943A;
wire g11171A;
wire I6631A;
wire g6064A;
wire g7230A;
wire g1648A;
wire g4952A;
wire g266A;
wire g6787A;
wire g8968A;
wire g10306A;
wire g11459A;
wire g538A;
wire g11458A;
wire g5739A;
wire g7496A;
wire g4986A;
wire g5187A;
wire g11010A;
wire g1741A;
wire g3999A;
wire g8175A;
wire g8722A;
wire g5590A;
wire g7471A;
wire g7891A;
wire g8651A;
wire g5479A;
wire g11599A;
wire g6684A;
wire g6745A;
wire g357A;
wire g6639A;
wire g3696A;
wire g4503A;
wire g6791A;
wire g8180A;
wire g1092A;
wire g4224A;
wire g5501A;
wire g8602A;
wire g8838A;
wire g10666A;
wire g309A;
wire g11158A;
wire g9602A;
wire g5704A;
wire g3879A;
wire g4617A;
wire g9868A;
wire g11295A;
wire g11144A;
wire g1540A;
wire g9718A;
wire g3434A;
wire g4987A;
wire g1270A;
wire g1065A;
wire g6098A;
wire g9582A;
wire g3533A;
wire g8104A;
wire g1733A;
wire g9415A;
wire g8377A;
wire g8499A;
wire g9664A;
wire g9413A;
wire g3584A;
wire g6162A;
wire g1508A;
wire g4991A;
wire g5846A;
wire g6362A;
wire g10685A;
wire g1153A;
wire g11023A;
wire g7598A;
wire g11224A;
wire g11571A;
wire g1520A;
wire g4959A;
wire g1633A;
wire g5626A;
wire g9920A;
wire g9940A;
wire g1086A;
wire g4876A;
wire g6730A;
wire g263A;
wire g9689A;
wire g10762A;
wire g1050A;
wire g6070A;
wire g9428A;
wire g1759A;
wire g9430A;
wire g8927A;
wire g7068A;
wire g7740A;
wire g8014A;
wire g11278A;
wire g5782A;
wire g4236A;
wire g11559A;
wire g9609A;
wire g11558A;
wire g6087A;
wire g10751A;
wire g10655A;
wire g10772A;
wire g8135A;
wire g11544A;
wire g5084A;
wire g8382A;
wire g10230A;
wire g7241A;
wire g3942A;
wire g10638A;
wire g4064A;
wire g1321A;
wire g9365A;
wire g9738A;
wire g9579A;
wire g9861A;
wire g11255A;
wire g11189A;
wire g10510A;
wire g2917A;
wire g11188A;
wire g9846A;
wire g1878A;
wire g7818A;
wire g11460A;
wire g11030A;
wire g841A;
wire g11093A;
wire g7478A;
wire g7893A;
wire g8653A;
wire g10442A;
wire g6535A;
wire g8102A;
wire g1490A;
wire g1494A;
wire I5085A;
wire g3912A;
wire g7186A;
wire g4489A;
wire g9662A;
wire g9418A;
wire g959A;
wire g11218A;
wire g1121A;
wire g10643A;
wire g10746A;
wire g7125A;
wire g7821A;
wire g6246A;
wire g8963A;
wire g7533A;
wire g10237A;
wire g7939A;
wire g8638A;
wire g8786A;
wire g10684A;
wire g11455A;
wire g8364A;
wire g2990A;
wire g9847A;
wire g7584A;
wire g5617A;
wire g5981A;
wire g5789A;
wire g4009A;
wire g11277A;
wire g6472A;
wire g6940A;
wire g6760A;
wire g7061A;
wire g11595A;
wire g5771A;
wire g8405A;
wire g8553A;
wire g4836A;
wire g5547A;
wire g4967A;
wire g342A;
wire g6671A;
wire g7200A;
wire g382A;
wire g7046A;
wire g999A;
wire g4229A;
wire g8389A;
wire g6430A;
wire g4993A;
wire g6247A;
wire g11170A;
wire g7145A;
wire g5738A;
wire g3998A;
wire g6741A;
wire g11167A;
wire g11194A;
wire g1333A;
wire g11589A;
wire g4431A;
wire g7536A;
wire g9585A;
wire g2957A;
wire g11588A;
wire g5690A;
wire g6883A;
wire g1068A;
wire g4837A;
wire g8641A;
wire g8791A;
wire g6217A;
wire g444A;
wire g11022A;
wire g4168A;
wire g5915A;
wire g511A;
wire g5110A;
wire g11254A;
wire g7567A;
wire g3273A;
wire g4392A;
wire g1592A;
wire g9856A;
wire g9411A;
wire g5002A;
wire g857A;
wire g11101A;
wire g11177A;
wire g11560A;
wire g8098A;
wire g3970A;
wire g4941A;
wire g366A;
wire g6662A;
wire g7935A;
wire g6067A;
wire g9740A;
wire g9863A;
wire g174A;
wire g170A;
wire g6758A;
wire g6994A;
wire g1589A;
wire g1007A;
wire g4252A;
wire g542A;
wire g11166A;
wire g7130A;
wire g5179A;
wire g11009A;
wire g7542A;
wire g5171A;
wire g11008A;
wire g1209A;
wire g3516A;
wire g7573A;
wire g3987A;
wire g491A;
wire g11555A;
wire g9734A;
wire g9569A;
wire g9857A;
wire g8728A;
wire g8730A;
wire g8185A;
wire g1610A;
wire g8385A;
wire g7902A;
wire g4073A;
wire g8070A;
wire g5731A;
wire g11238A;
wire g1125A;
wire g8308A;
wire g8470A;
wire g5489A;
wire g3991A;
wire g166A;
wire g7823A;
wire g4069A;
wire g1317A;
wire g11176A;
wire g837A;
wire g11092A;
wire g330A;
wire g11154A;
wire g7A;
wire g9608A;
wire g11637A;
wire g2091A;
wire g8406A;
wire g5254A;
wire g8612A;
wire g9588A;
wire g8742A;
wire g8801A;
wire g7063A;
wire g10303A;
wire g1486A;
wire g5009A;
wire g9665A;
wire g8748A;
wire g11215A;
wire g10750A;
wire g3818A;
wire g5769A;
wire g6673A;
wire g1255A;
wire g7720A;
wire g4609A;
wire g7547A;
wire g7971A;
wire g11288A;
wire g7599A;
wire g6058A;
wire g4106A;
wire g6743A;
wire g6890A;
wire g7269A;
wire g7549A;
wire g8169A;
wire g11304A;
wire g9924A;
wire g9944A;
wire g7592A;
wire g8718A;
wire g8616A;
wire g9316A;
wire g7625A;
wire g8644A;
wire g8793A;
wire g2940A;
wire g11624A;
wire g2947A;
wire g10949A;
wire g3563A;
wire g2223A;
wire g10948A;
wire g7846A;
wire g8246A;
wire g5788A;
wire g4008A;
wire g9596A;
wire g5249A;
wire g11585A;
wire g4972A;
wire g11554A;
wire g7096A;
wire g10673A;
wire g2493A;
wire g4806A;
wire g9915A;
wire g9936A;
wire g1660A;
wire g2910A;
wire g9317A;
wire g10853A;
wire g10933A;
wire g8177A;
wire g8388A;
wire g1117A;
wire g7141A;
wire g10508A;
wire g4230A;
wire g10634A;
wire g9192A;
wire g9601A;
wire g6326A;
wire g700A;
wire g7710A;
wire g7375A;
wire g8028A;
wire g5640A;
wire g5031A;
wire g4550A;
wire g7879A;
wire g7962A;
wire g9597A;
wire g631A;
wire g5005A;
wire g6423A;
wire g8108A;
wire g3322A;
wire g5911A;
wire g9916A;
wire g9937A;
wire g9704A;
wire g9747A;
wire g9840A;
wire g10723A;
wire g8217A;
wire g5209A;
wire g11013A;
wire g9390A;
wire g11214A;
wire g6327A;
wire g1149A;
wire g5796A;
wire g5473A;
wire g5038A;
wire g6346A;
wire g6633A;
wire g5119A;
wire g11005A;
wire g8365A;
wire g7558A;
wire g4481A;
wire g4097A;
wire g7588A;
wire g4497A;
wire g9922A;
wire g9942A;
wire g6696A;
wire g5118A;
wire g1850A;
wire g10665A;
wire g10731A;
wire g8552A;
wire g8827A;
wire g5540A;
wire g1403A;
wire g4960A;
wire g8615A;
wire g8846A;
wire g5983A;
wire g182A;
wire g6240A;
wire g7931A;
wire g853A;
wire g11100A;
wire g11235A;
wire g5199A;
wire g6316A;
wire g7515A;
wire g5781A;
wire g7742A;
wire g8018A;
wire g2950A;
wire g5510A;
wire g6347A;
wire g962A;
wire g9357A;
wire g11407A;
wire g10743A;
wire g5259A;
wire g5694A;
wire g10769A;
wire g11584A;
wire g4932A;
wire g10649A;
wire g10768A;
wire g4068A;
wire g6317A;
wire g4276A;
wire g5215A;
wire g6775A;
wire g10662A;
wire g8101A;
wire g3204A;
wire g5318A;
wire g5825A;
wire g7457A;
wire g7884A;
wire g1292A;
wire g3974A;
wire g9929A;
wire g9949A;
wire g10778A;
wire g7524A;
wire g6079A;
wire g7235A;
wire g9603A;
wire g9726A;
wire g9850A;
wire g7988A;
wire g5228A;
wire g5587A;
wire g5934A;
wire g8168A;
wire g9583A;
wire g10672A;
wire g8627A;
wire g635A;
wire g8309A;
wire g10449A;
wire g11273A;
wire g8734A;
wire g5913A;
wire g4572A;
wire g6363A;
wire g11463A;
wire g718A;
wire g8074A;
wire g1166A;
wire g8383A;
wire g8474A;
wire g11234A;
wire g4483A;
wire g11491A;
wire g5097A;
wire g5726A;
wire g5497A;
wire g7933A;
wire g9A;
wire g9617A;
wire g9873A;
wire g9906A;
wire g5196A;
wire g11012A;
wire g7050A;
wire g10849A;
wire g10971A;
wire g8400A;
wire g1169A;
wire g4345A;
wire g9925A;
wire g9945A;
wire g5028A;
wire g7271A;
wire g9709A;
wire g1003A;
wire g4223A;
wire g10497A;
wire g10716A;
wire g11247A;
wire g6661A;
wire g11173A;
wire g6075A;
wire g7367A;
wire g8023A;
wire g9888A;
wire g9907A;
wire g10582A;
wire g5746A;
wire g9950A;
wire g9959A;
wire g7674A;
wire g9690A;
wire g5703A;
wire g360A;
wire g4522A;
wire g4115A;
wire g7075A;
wire g10627A;
wire g4047A;
wire g2944A;
wire g6646A;
wire g7132A;
wire g11029A;
wire g7572A;
wire g8127A;
wire g7209A;
wire g11028A;
wire g10742A;
wire g8880A;
wire g10681A;
wire g9663A;
wire g5349A;
wire g8732A;
wire g3807A;
wire g3860A;
wire g5848A;
wire g8411A;
wire g8508A;
wire g8072A;
wire g5699A;
wire g11240A;
wire g6105A;
wire g6616A;
wire g10690A;
wire g7582A;
wire g9590A;
wire g4128A;
wire g6404A;
wire g6647A;
wire g10504A;
wire g9657A;
wire g4542A;
wire g1163A;
wire g5524A;
wire g9899A;
wire g7736A;
wire g10626A;
wire g6320A;
wire g7623A;
wire g10299A;
wire g7889A;
wire g10298A;
wire g8413A;
wire g3979A;
wire g1848A;
wire g5211A;
wire g4512A;
wire g7722A;
wire g9714A;
wire g9522A;
wire g9844A;
wire g1141A;
wire g5993A;
wire g5026A;
wire g8705A;
wire g10737A;
wire g10232A;
wire g6771A;
wire g5170A;
wire g8117A;
wire g9956A;
wire g9966A;
wire g5280A;
wire g7139A;
wire g11099A;
wire g6892A;
wire g9705A;
wire g10512A;
wire g849A;
wire g11098A;
wire g8628A;
wire g5544A;
wire g11272A;
wire g1621A;
wire g5483A;
wire g9928A;
wire g9948A;
wire g4063A;
wire g11462A;
wire g6738A;
wire g7593A;
wire g11032A;
wire g10445A;
wire g8882A;
wire g10316A;
wire g5756A;
wire g1023A;
wire g4720A;
wire g9409A;
wire g8929A;
wire g6876A;
wire g4989A;
wire g9737A;
wire g9836A;
wire g6061A;
wire g8268A;
wire g6465A;
wire g1466A;
wire g5003A;
wire g9957A;
wire g9967A;
wire g5145A;
wire g4971A;
wire g10753A;
wire g5695A;
wire g7613A;
wire g10736A;
wire g11220A;
wire g7444A;
wire g4670A;
wire g4253A;
wire g7960A;
wire g8163A;
wire g10764A;
wire g5757A;
wire g7385A;
wire g8032A;
wire g2988A;
wire g11591A;
wire g7583A;
wire g321A;
wire g11147A;
wire g5522A;
wire g1394A;
wire g9697A;
wire g9751A;
wire g9837A;
wire g9620A;
wire g327A;
wire g11151A;
wire g11172A;
wire g7885A;
wire g5595A;
wire g5537A;
wire g9708A;
wire g9516A;
wire g9842A;
wire g4141A;
wire g4341A;
wire g7679A;
wire g7378A;
wire g5612A;
wire g7135A;
wire g10970A;
wire g11025A;
wire g9730A;
wire g9854A;
wire g7182A;
wire g9921A;
wire g9941A;
wire g6194A;
wire g1651A;
wire g4962A;
wire g4358A;
wire g4803A;
wire g8549A;
wire g8683A;
wire g1113A;
wire g5224A;
wire g8778A;
wire g11281A;
wire g318A;
wire g11146A;
wire g2948A;
wire g3904A;
wire g8075A;
wire g9723A;
wire g9829A;
wire g7184A;
wire g11246A;
wire g5837A;
wire g6350A;
wire g2555A;
wire g5902A;
wire g1765A;
wire g6438A;
wire g5512A;
wire g5090A;
wire g7719A;
wire g3695A;
wire g7587A;
wire g9610A;
wire g3536A;
wire g8881A;
wire g4559A;
wire g10549A;
wire g10561A;
wire g5698A;
wire g11226A;
wire g10295A;
wire g5260A;
wire g10680A;
wire g1853A;
wire g11538A;
wire g11551A;
wire g9849A;
wire g5279A;
wire g8404A;
wire g5720A;
wire g11318A;
wire g11297A;
wire g9898A;
wire g9510A;
wire g7297A;
wire g7963A;
wire g9759A;
wire g9803A;
wire g11338A;
wire g8435A;
wire g6124A;
wire I5600A;
wire g11257A;
wire g11256A;
wire g3107A;
wire g2167A;
wire I14866A;
wire g4997A;
wire g10291A;
wire g6122A;
wire g9509A;
wire g5227A;
wire I15054A;
wire g11269A;
wire g5555A;
wire g11268A;
wire g11335A;
wire g8249A;
wire g9882A;
wire I15210A;
wire g2102A;
wire g2099A;
wire g2096A;
wire g2088A;
wire I5805A;
wire g11443A;
wire g8431A;
wire g8286A;
wire g7290A;
wire g8287A;
wire g7301A;
wire g8259A;
wire g11334A;
wire g10805A;
wire I15214A;
wire I15215A;
wire g11265A;
wire g8322A;
wire g8433A;
wire g8248A;
wire g8154A;
wire g2405A;
wire g2389A;
wire g2380A;
wire g2372A;
wire I6351A;
wire I16427A;
wire g7303A;
wire g2862A;
wire g2515A;
wire g4052A;
wire I14858A;
wire g11264A;
wire I15209A;
wire g1570A;
wire g2528A;
wire g2522A;
wire g9515A;
wire g7294A;
wire g3118A;
wire g2180A;
wire I5571A;
wire I5599A;
wire g2514A;
wire g11327A;
wire I5629A;
wire I5363A;
wire g2315A;
wire g8159A;
wire g11326A;
wire I16148A;
wire I16149A;
wire g10521A;
wire g7292A;
wire g8417A;
wire I14855A;
wire g9878A;
wire I15205A;
wire I15051A;
wire g8823A;
wire g8148A;
wire g2863A;
wire g2516A;
wire g7299A;
wire g9511A;
wire g9654A;
wire I15224A;
wire I15225A;
wire g8253A;
wire I15171A;
wire I15172A;
wire I15204A;
wire g10472A;
wire g10470A;
wire g10468A;
wire g10467A;
wire g10386A;
wire g10384A;
wire g10476A;
wire g10474A;
wire g8158A;
wire g11331A;
wire g7295A;
wire g8284A;
wire g1393A;
wire I5357A;
wire g9758A;
wire I5626A;
wire g7298A;
wire g8282A;
wire I15057A;
wire I15219A;
wire I15220A;
wire I14862A;
wire g2521A;
wire g9591A;
wire g9757A;
wire g11261A;
wire g9815A;
wire I14835A;
wire g126A;
wire g10479A;
wire g10478A;
wire g10477A;
wire g10475A;
wire I16161A;
wire g2353A;
wire I5804A;
wire g7291A;
wire I15199A;
wire g11330A;
wire g8153A;
wire g9881A;
wire g11259A;
wire g11258A;
wire g9426A;
wire g9423A;
wire g11337A;
wire g8262A;
wire g8285A;
wire I5570A;
wire g2499A;
wire g11336A;
wire g7293A;
wire g9388A;
wire g11260A;
wire g10807A;
wire g8288A;
wire g10394A;
wire g10392A;
wire g10482A;
wire g10481A;
wire I16160A;
wire g9589A;
wire g11270A;
wire g11267A;
wire g1959A;
wire g9667A;
wire I14827A;
wire g9391A;
wire I5358A;
wire g2309A;
wire g11266A;
wire g8429A;
wire g8281A;
wire g9876A;
wire I15177A;
wire g5186A;
wire I6350A;
wire g1527A;
wire g8162A;
wire I14779A;
wire I5351A;
wire I5352A;
wire g2305A;
wire I15176A;
wire g9879A;
wire g8283A;
wire g11333A;
wire g10562A;
wire g9606A;
wire I14822A;
wire g9880A;
wire I15200A;
wire g8428A;
wire g8430A;
wire g8247A;
wire I5576A;
wire g4476A;
wire I5649A;
wire g2538A;
wire g11329A;
wire g11328A;
wire g9605A;
wire g9363A;
wire g7300A;
wire I14831A;
wire g8263A;
wire g11263A;
wire g5780A;
wire g11332A;
wire I15048A;
wire g9647A;
wire I14602A;
wire I15033A;
wire g2445A;
wire g2437A;
wire g2433A;
wire g2419A;
wire g11325A;
wire I5366A;
wire g9506A;
wire g8161A;
wire g2316A;
wire g4675A;
wire g8434A;
wire g11262A;
wire g9387A;
wire I15045A;
wire g11324A;
wire g2501A;
wire g9877A;
wire g10529A;
wire g8432A;
wire g9874A;
wire g8157A;
wire g6899A;
wire g9646A;
wire g7302A;
wire g2111A;
wire g2109A;
wire g2106A;
wire g2104A;
wire g7296A;
wire I5612A;
wire I5613A;
wire I5591A;
wire I5593A;
wire g8839A;
wire g8970A;
wire I10519A;
wire I11278A;
wire I11279A;
wire g3978A;
wire I5263A;
wire I5264A;
wire g4278A;
wire I8640A;
wire g2943A;
wire I6760A;
wire I6761A;
wire g11418A;
wire g11416A;
wire I17400A;
wire I5449A;
wire I5450A;
wire I16058A;
wire I16060A;
wire g2938A;
wire I6746A;
wire I11973A;
wire I11975A;
wire I12136A;
wire I11935A;
wire I11937A;
wire I6167A;
wire I6168A;
wire g2959A;
wire g2120A;
wire g2115A;
wire I5878A;
wire I5619A;
wire I5620A;
wire g5552A;
wire I6467A;
wire I6468A;
wire g4672A;
wire I8795A;
wire I8796A;
wire I15891A;
wire I15892A;
wire I5611A;
wire g8738A;
wire I6714A;
wire I6716A;
wire g3460A;
wire I7683A;
wire I7685A;
wire I12106A;
wire I12108A;
wire I6747A;
wire I5230A;
wire I5231A;
wire g2236A;
wire I12075A;
wire I12076A;
wire I15870A;
wire I16065A;
wire I16067A;
wire I7562A;
wire I13529A;
wire I13531A;
wire I8797A;
wire I17584A;
wire I11936A;
wire I15256A;
wire I15257A;
wire I13505A;
wire I13506A;
wire g8502A;
wire g8501A;
wire g8824A;
wire I6186A;
wire I17504A;
wire I17505A;
wire g11496A;
wire I15999A;
wire I16001A;
wire g2215A;
wire I6124A;
wire I6125A;
wire I11907A;
wire I11909A;
wire I12038A;
wire I12040A;
wire I13907A;
wire I13909A;
wire I6771A;
wire I6772A;
wire I11908A;
wire I16008A;
wire I16009A;
wire I13908A;
wire I7034A;
wire I7035A;
wire I8650A;
wire I9947A;
wire I9948A;
wire g10428A;
wire I16066A;
wire I6144A;
wire I6145A;
wire I11241A;
wire I11242A;
wire I15993A;
wire I15994A;
wire I6187A;
wire g6027A;
wire I5500A;
wire I11974A;
wire I12060A;
wire I12062A;
wire I8771A;
wire I8772A;
wire I5184A;
wire I13293A;
wire I6199A;
wire I6200A;
wire I13265A;
wire I5023A;
wire I5024A;
wire I7863A;
wire I13991A;
wire I13992A;
wire I13660A;
wire I13661A;
wire I6143A;
wire I13990A;
wire I11508A;
wire I11510A;
wire g5034A;
wire I5229A;
wire I12045A;
wire I12047A;
wire I10769A;
wire I10771A;
wire I16045A;
wire I16046A;
wire I12061A;
wire I5104A;
wire I13530A;
wire I6447A;
wire I4954A;
wire I4956A;
wire g3530A;
wire I8479A;
wire I8481A;
wire I8739A;
wire I8740A;
wire I6879A;
wire I6880A;
wire I15430A;
wire I15431A;
wire I12019A;
wire I12020A;
wire I16331A;
wire I16332A;
wire I16467A;
wire I16469A;
wire I5013A;
wire I5014A;
wire I13521A;
wire I13523A;
wire I16037A;
wire I16039A;
wire I16468A;
wire I12046A;
wire I16038A;
wire g4374A;
wire I8676A;
wire I12113A;
wire g4616A;
wire I8761A;
wire I15992A;
wire I5034A;
wire I5036A;
wire g8843A;
wire I14263A;
wire I13249A;
wire I13250A;
wire I5135A;
wire I5485A;
wire I5486A;
wire I7033A;
wire I15441A;
wire I15443A;
wire I6166A;
wire g4267A;
wire I8624A;
wire I16015A;
wire I8677A;
wire g4234A;
wire I8575A;
wire I8576A;
wire g9204A;
wire I14612A;
wire I14613A;
wire g4601A;
wire I8715A;
wire I8716A;
wire I6715A;
wire I13514A;
wire I13515A;
wire I12002A;
wire I12003A;
wire I5127A;
wire I5128A;
wire g2177A;
wire I8577A;
wire g11414A;
wire I17393A;
wire I17395A;
wire I11280A;
wire I5265A;
wire I6988A;
wire I6989A;
wire I13272A;
wire I13274A;
wire I10507A;
wire I5164A;
wire I14443A;
wire I14444A;
wire I9557A;
wire I9559A;
wire I5592A;
wire I13077A;
wire I13078A;
wire I8717A;
wire I5295A;
wire I5296A;
wire I8625A;
wire I8626A;
wire I4911A;
wire I4912A;
wire I16000A;
wire I5371A;
wire I5185A;
wire I5186A;
wire I5675A;
wire g4218A;
wire I8543A;
wire I8544A;
wire I10520A;
wire I10521A;
wire I5297A;
wire I13537A;
wire I13283A;
wire g4749A;
wire I11980A;
wire I11982A;
wire g4873A;
wire I8513A;
wire I8514A;
wire I13089A;
wire I13091A;
wire I6126A;
wire g10302A;
wire I15906A;
wire I15908A;
wire I8763A;
wire g8506A;
wire g8825A;
wire I16007A;
wire g2107A;
wire g2105A;
wire I5865A;
wire I5604A;
wire I5517A;
wire I5518A;
wire I6109A;
wire I6111A;
wire I4929A;
wire I4930A;
wire I13522A;
wire I10770A;
wire I5538A;
wire I5539A;
wire g11415A;
wire I17394A;
wire I13552A;
wire I13553A;
wire I8642A;
wire I17296A;
wire I17297A;
wire I14278A;
wire I14279A;
wire I4910A;
wire I6792A;
wire I6794A;
wire I5484A;
wire I15442A;
wire I10931A;
wire I10932A;
wire I8779A;
wire I8780A;
wire g2354A;
wire g10043A;
wire g10153A;
wire I15615A;
wire I17281A;
wire I5468A;
wire I5470A;
wire I11509A;
wire I5025A;
wire I14270A;
wire I14272A;
wire I6208A;
wire I6209A;
wire I17288A;
wire I17290A;
wire I7563A;
wire I7564A;
wire I5005A;
wire I5006A;
wire I12126A;
wire I12128A;
wire I5105A;
wire I6322A;
wire I6323A;
wire I12093A;
wire I12094A;
wire g2776A;
wire I6664A;
wire I6666A;
wire I6762A;
wire g3623A;
wire I5373A;
wire I8527A;
wire I8529A;
wire I5282A;
wire I5283A;
wire I7223A;
wire I7224A;
wire I5007A;
wire I5459A;
wire I17295A;
wire I5015A;
wire I14264A;
wire I14265A;
wire I16072A;
wire I16073A;
wire g3205A;
wire I8652A;
wire I9558A;
wire I5202A;
wire I5203A;
wire I6806A;
wire I6807A;
wire I6469A;
wire I12143A;
wire I12145A;
wire I12127A;
wire I13300A;
wire I13302A;
wire I5502A;
wire I9574A;
wire I6448A;
wire I6449A;
wire I8669A;
wire I8670A;
wire I15451A;
wire I15453A;
wire I7875A;
wire I7876A;
wire I14202A;
wire I14203A;
wire g10149A;
wire g10144A;
wire I15607A;
wire I5324A;
wire I5325A;
wire I8738A;
wire g10434A;
wire g5859A;
wire I8604A;
wire I8606A;
wire I12085A;
wire I12087A;
wire I13248A;
wire I4979A;
wire I4980A;
wire I12067A;
wire I12069A;
wire g8942A;
wire I12068A;
wire I17503A;
wire I7877A;
wire I5165A;
wire I6287A;
wire I6289A;
wire I6777A;
wire I8562A;
wire I8563A;
wire I15890A;
wire g8006A;
wire I13090A;
wire I17460A;
wire I17461A;
wire g11474A;
wire I13513A;
wire I4986A;
wire I4987A;
wire I5204A;
wire I13504A;
wire I6207A;
wire I12086A;
wire I8545A;
wire I8178A;
wire I8180A;
wire I8589A;
wire I8591A;
wire I10930A;
wire I17402A;
wire I13294A;
wire I13295A;
wire I12144A;
wire g8757A;
wire g2961A;
wire I14209A;
wire I14211A;
wire I8515A;
wire I5316A;
wire I5317A;
wire I9946A;
wire g4613A;
wire I8750A;
wire I5605A;
wire I14204A;
wire I16051A;
wire g10360A;
wire g6037A;
wire I13858A;
wire I13859A;
wire I15872A;
wire g4879A;
wire I8528A;
wire I13901A;
wire I13902A;
wire g8542A;
wire I6836A;
wire I6838A;
wire I17305A;
wire I17307A;
wire g4538A;
wire I15452A;
wire I13857A;
wire I13765A;
wire I8671A;
wire I16044A;
wire g10363A;
wire g5360A;
wire I5106A;
wire g4677A;
wire I8803A;
wire I8804A;
wire I16016A;
wire I16017A;
wire I17485A;
wire I17487A;
wire I4995A;
wire I12092A;
wire I8678A;
wire I5126A;
wire I5372A;
wire I17306A;
wire I11995A;
wire I7225A;
wire I11261A;
wire g8545A;
wire I6110A;
wire I4941A;
wire I4942A;
wire I15899A;
wire I15900A;
wire g5527A;
wire g5350A;
wire I16079A;
wire I16081A;
wire I8641A;
wire I6176A;
wire I6178A;
wire I12074A;
wire I5451A;
wire I7322A;
wire I7323A;
wire I6288A;
wire I8179A;
wire I6805A;
wire I17486A;
wire I4928A;
wire I16330A;
wire I9575A;
wire I13886A;
wire I13887A;
wire I8787A;
wire I8788A;
wire I5315A;
wire g10285A;
wire I13867A;
wire I13869A;
wire I13868A;
wire I13258A;
wire I13259A;
wire g3261A;
wire I16074A;
wire I5136A;
wire I5137A;
wire I5460A;
wire I5461A;
wire I8605A;
wire I6770A;
wire I17401A;
wire g11449A;
wire g11448A;
wire g10231A;
wire I15716A;
wire I15717A;
wire I14210A;
wire I17567A;
wire I17569A;
wire I13876A;
wire I13878A;
wire I5606A;
wire I14442A;
wire I11996A;
wire I11997A;
wire I14277A;
wire I17568A;
wire I7321A;
wire I6990A;
wire g8847A;
wire I9006A;
wire I4985A;
wire I8651A;
wire I13544A;
wire I13545A;
wire I13894A;
wire I13895A;
wire I6136A;
wire I6138A;
wire I13076A;
wire g2205A;
wire I13260A;
wire I5501A;
wire I17586A;
wire I13900A;
wire I6201A;
wire g8826A;
wire I14216A;
wire I14217A;
wire I9007A;
wire I13559A;
wire I13561A;
wire g10229A;
wire I17492A;
wire I17493A;
wire I12214A;
wire I12215A;
wire I11262A;
wire I11263A;
wire I6225A;
wire I6226A;
wire I13307A;
wire I13309A;
wire I5676A;
wire I5677A;
wire I6826A;
wire I6827A;
wire g8190A;
wire I13308A;
wire I5879A;
wire I5880A;
wire g2792A;
wire g3061A;
wire I17585A;
wire I6881A;
wire I12138A;
wire g4605A;
wire I8728A;
wire I8729A;
wire I15871A;
wire I5866A;
wire I5867A;
wire I6793A;
wire I6487A;
wire I16080A;
wire I13893A;
wire I12115A;
wire I6748A;
wire I6224A;
wire I8805A;
wire I15878A;
wire I15880A;
wire I16030A;
wire I16031A;
wire I14271A;
wire I13267A;
wire I15616A;
wire I15617A;
wire I4964A;
wire I4966A;
wire I8752A;
wire I15432A;
wire g10438A;
wire g6032A;
wire g3011A;
wire I8480A;
wire I16086A;
wire I16087A;
wire g3734A;
wire I14218A;
wire I4955A;
wire g4639A;
wire I8786A;
wire g10480A;
wire I11914A;
wire I11915A;
wire g4619A;
wire I8770A;
wire I5516A;
wire g8541A;
wire I6188A;
wire I5891A;
wire I5892A;
wire I13766A;
wire I13767A;
wire I15258A;
wire I13266A;
wire I6825A;
wire I17283A;
wire g5277A;
wire I5035A;
wire g10359A;
wire I15879A;
wire I12114A;
wire I12107A;
wire g2500A;
wire g10430A;
wire g5999A;
wire I13285A;
wire I13877A;
wire I5893A;
wire g2795A;
wire I13560A;
wire g4259A;
wire I5166A;
wire I14614A;
wire I4965A;
wire I4943A;
wire I16023A;
wire I16059A;
wire g8737A;
wire I9576A;
wire I16052A;
wire I16053A;
wire I12004A;
wire g5573A;
wire I6837A;
wire I8730A;
wire I4978A;
wire I6177A;
wire I17051A;
wire I7864A;
wire I7865A;
wire I6665A;
wire I12216A;
wire I13554A;
wire I13284A;
wire I6137A;
wire I5529A;
wire I5530A;
wire I17282A;
wire I5618A;
wire I8662A;
wire I8664A;
wire I11916A;
wire g7717A;
wire I4971A;
wire I4972A;
wire I13273A;
wire I10509A;
wire I10508A;
wire I6778A;
wire I6779A;
wire I5469A;
wire g4251A;
wire I13546A;
wire I4996A;
wire I4997A;
wire I13539A;
wire I16032A;
wire I5323A;
wire I13538A;
wire I5540A;
wire I8778A;
wire g4286A;
wire I17052A;
wire I17053A;
wire I15898A;
wire g7978A;
wire g4227A;
wire I8561A;
wire I8762A;
wire I8751A;
wire I15907A;
wire I4973A;
wire I16024A;
wire I16025A;
wire g4455A;
wire I5341A;
wire I5342A;
wire I12137A;
wire I16088A;
wire g10483A;
wire I17289A;
wire g4630A;
wire I15609A;
wire I15608A;
wire g10436A;
wire g6023A;
wire I17459A;
wire I13301A;
wire I11981A;
wire I8663A;
wire I15718A;
wire I5284A;
wire g4607A;
wire g8840A;
wire g10441A;
wire g5345A;
wire g10432A;
wire g5938A;
wire I12021A;
wire I6489A;
wire I5528A;
wire I13659A;
wire I5343A;
wire I12039A;
wire I9008A;
wire I6488A;
wire I13888A;
wire I17494A;
wire I7684A;
wire g3221A;
wire I6324A;
wire I8590A;
wire I11243A;
wire g1737A;
wire g10324A;
wire g10239A;
wire g4974A;
wire g10322A;
wire g1736A;
wire g1955A;
wire g1956A;
wire g113A;
wire g1360A;
wire g1217A;
wire g755A;
wire g875A;
wire g1356A;
wire g874A;
wire FE_OFN370_g4525B;
wire FE_OFN369_g4525B;
wire FE_OFN368_g4525B;
wire FE_OFN367_g3521B;
wire FE_OFN366_g3521B;
wire FE_OFN365_g5361B;
wire FE_OFN364_g3015B;
wire FE_OFN363_I5565B;
wire FE_OFN362_g4525B;
wire FE_OFN360_g4525B;
wire FE_OFN359_g18B;
wire FE_OFN358_g3521B;
wire FE_OFN357_g3521B;
wire FE_OFN356_g5361B;
wire FE_OFN354_g5361B;
wire FE_OFN353_g5117B;
wire FE_OFN352_g109B;
wire FE_OFN351_g3913B;
wire FE_OFN350_g3121B;
wire FE_OFN349_I6424B;
wire FE_OFN348_g3015B;
wire FE_OFN347_g3914B;
wire FE_OFN346_g4381B;
wire FE_OFN345_g3015B;
wire FE_OFN344_g3586B;
wire FE_OFN343_I5565B;
wire FE_OFN340_I5565B;
wire FE_OFN339_g4525B;
wire FE_OFN337_g4525B;
wire FE_OFN336_g1690B;
wire FE_OFN335_g4737B;
wire FE_OFN334_g7045B;
wire FE_OFN333_g4294B;
wire FE_OFN332_g8748B;
wire FE_OFN331_g8696B;
wire FE_OFN330_g7638B;
wire FE_OFN329_g8763B;
wire FE_OFN328_g8709B;
wire FE_OFN325_g18B;
wire FE_OFN324_g18B;
wire FE_OFN322_g4449B;
wire FE_OFN321_g5261B;
wire FE_OFN320_g5361B;
wire FE_OFN319_g5361B;
wire FE_OFN318_g5361B;
wire FE_OFN316_g5361B;
wire FE_OFN315_g5117B;
wire FE_OFN312_g5117B;
wire FE_OFN310_g4336B;
wire FE_OFN308_I6424B;
wire FE_OFN307_g4010B;
wire FE_OFN306_g5128B;
wire FE_OFN305_g5151B;
wire FE_OFN304_g5151B;
wire FE_OFN303_g4678B;
wire FE_OFN302_g3913B;
wire FE_OFN300_g4002B;
wire FE_OFN299_g4457B;
wire FE_OFN298_g3015B;
wire FE_OFN297_g3015B;
wire FE_OFN296_g3914B;
wire FE_OFN294_g3914B;
wire FE_OFN293_g3015B;
wire FE_OFN292_g3015B;
wire FE_OFN291_g4880B;
wire FE_OFN290_g4880B;
wire FE_OFN289_g4679B;
wire FE_OFN288_g4263B;
wire FE_OFN287_g3586B;
wire FE_OFN284_g3586B;
wire FE_OFN283_I8869B;
wire FE_OFN282_g6165B;
wire FE_OFN281_g2216B;
wire FE_OFN280_g9536B;
wire FE_OFN279_g11157B;
wire FE_OFN278_g10927B;
wire FE_OFN277_g48B;
wire FE_OFN276_g48B;
wire FE_OFN275_g48B;
wire FE_OFN273_g85B;
wire FE_OFN271_g85B;
wire FE_OFN269_g109B;
wire FE_OFN267_g109B;
wire FE_OFN266_g18B;
wire FE_OFN260_g18B;
wire FE_OFN254_g461B;
wire FE_OFN253_g1786B;
wire FE_OFN252_g1791B;
wire FE_OFN251_g1801B;
wire FE_OFN250_g471B;
wire FE_OFN248_g466B;
wire FE_OFN247_g1771B;
wire FE_OFN245_g1690B;
wire FE_OFN241_g1690B;
wire FE_OFN240_g1110B;
wire FE_OFN239_g1796B;
wire FE_OFN238_g1781B;
wire FE_OFN237_g1806B;
wire FE_OFN236_g1776B;
wire FE_OFN235_g2024B;
wire FE_OFN234_g2024B;
wire FE_OFN233_I5565B;
wire FE_OFN230_I5565B;
wire FE_OFN229_g3880B;
wire FE_OFN227_g3880B;
wire FE_OFN226_g3880B;
wire FE_OFN225_g2276B;
wire FE_OFN224_g2276B;
wire FE_OFN223_g4401B;
wire FE_OFN221_g3440B;
wire FE_OFN219_g5557B;
wire FE_OFN218_g5557B;
wire FE_OFN217_g5013B;
wire FE_OFN213_g6003B;
wire FE_OFN211_g7246B;
wire FE_OFN210_g7246B;
wire FE_OFN209_g6863B;
wire FE_OFN207_g6863B;
wire FE_OFN206_g6863B;
wire FE_OFN204_g3664B;
wire FE_OFN200_g4921B;
wire FE_OFN199_g7697B;
wire FE_OFN198_g7697B;
wire FE_OFN196_g7697B;
wire FE_OFN195_g6488B;
wire FE_OFN192_g6488B;
wire FE_OFN191_g6488B;
wire FE_OFN189_g7638B;
wire FE_OFN187_g7638B;
wire FE_OFN184_I7048B;
wire FE_OFN180_g5354B;
wire FE_OFN179_g5354B;
wire FE_OFN178_g5354B;
wire FE_OFN177_g5919B;
wire FE_OFN176_g5151B;
wire FE_OFN168_g5361B;
wire FE_OFN166_g5361B;
wire FE_OFN164_g5361B;
wire FE_OFN161_g5361B;
wire FE_OFN160_I6424B;
wire FE_OFN155_g3121B;
wire FE_OFN154_g4640B;
wire FE_OFN153_g4640B;
wire FE_OFN147_g4682B;
wire FE_OFN146_g4682B;
wire FE_OFN144_g4682B;
wire FE_OFN142_g4682B;
wire FE_OFN141_g3829B;
wire FE_OFN137_g3829B;
wire FE_OFN136_g3863B;
wire FE_OFN134_g3863B;
wire FE_OFN133_g3015B;
wire FE_OFN132_g3015B;
wire FE_OFN131_g3015B;
wire FE_OFN119_g3015B;
wire FE_OFN118_g4807B;
wire FE_OFN117_g4807B;
wire FE_OFN116_g4807B;
wire FE_OFN115_g4807B;
wire FE_OFN113_g3914B;
wire FE_OFN111_g3914B;
wire FE_OFN110_g3586B;
wire FE_OFN103_g3586B;
wire FE_OFN102_g3586B;
wire FE_OFN100_g4421B;
wire FE_OFN99_g4421B;
wire FE_OFN97_I8869B;
wire FE_OFN96_g2169B;
wire FE_OFN95_g2216B;
wire FE_OFN93_g2216B;
wire FE_OFN92_g2216B;
wire FE_OFN91_g2172B;
wire FE_OFN90_I11360B;
wire FE_OFN89_I11360B;
wire FE_OFN88_g2178B;
wire FE_OFN87_g2176B;
wire FE_OFN86_g2176B;
wire FE_OFN85_g2176B;
wire FE_OFN84_g2176B;
wire FE_OFN83_g2176B;
wire FE_OFN82_g2176B;
wire FE_OFN81_g2176B;
wire FE_OFN80_g2175B;
wire FE_OFN79_g8700B;
wire FE_OFN76_g8700B;
wire FE_OFN73_g8858B;
wire FE_OFN72_g9292B;
wire FE_OFN71_g9292B;
wire FE_OFN70_g9490B;
wire FE_OFN69_g9392B;
wire FE_OFN68_g9392B;
wire FE_OFN67_g9367B;
wire FE_OFN64_g9536B;
wire FE_OFN63_g9474B;
wire FE_OFN62_g9274B;
wire FE_OFN61_g9624B;
wire FE_OFN60_g9624B;
wire FE_OFN59_g9432B;
wire FE_OFN57_g9432B;
wire FE_OFN56_g9052B;
wire FE_OFN54_g9052B;
wire FE_OFN53_g9173B;
wire FE_OFN52_g9173B;
wire FE_OFN51_g9111B;
wire FE_OFN50_g9030B;
wire FE_OFN49_g9030B;
wire FE_OFN48_g9151B;
wire FE_OFN47_g9151B;
wire FE_OFN46_g9125B;
wire FE_OFN45_g9125B;
wire FE_OFN44_g9125B;
wire FE_OFN42_g9205B;
wire FE_OFN40_g9240B;
wire FE_OFN39_g9223B;
wire FE_OFN35_g9785B;
wire FE_OFN34_g9785B;
wire FE_OFN33_g9454B;
wire FE_OFN32_g9454B;
wire FE_OFN27_g11519B;
wire FE_OFN21_g10702B;
wire FE_OFN20_g10702B;
wire FE_OFN18_g10702B;
wire FE_OFN17_g10702B;
wire FE_OFN15_g10702B;
wire FE_OFN14_g10702B;
wire FE_OFN13_g10702B;
wire FE_OFN10_g10702B;
wire FE_OFN9_g10702B;
wire FE_OFN8_g10702B;
wire FE_OFN7_g10702B;
wire FE_OFN4_g10950B;
wire FE_OFN3_g10950B;
wire FE_OFN0_g10950B;
wire g4500B;
wire g5529B;
wire g9968B;
wire g4682B;
wire g1707B;
wire g2299B;
wire g9291B;
wire g2807B;
wire I7048B;
wire g4130B;
wire g5024B;
wire g4338B;
wire g11596B;
wire g8147B;
wire g6551B;
wire g10865B;
wire g650B;
wire g1981B;
wire g8054B;
wire g3982B;
wire g9974B;
wire g1216B;
wire g546B;
wire g798B;
wire g3629B;
wire g7709B;
wire g8465B;
wire g8617B;
wire g4940B;
wire g4640B;
wire g135B;
wire g2078B;
wire g4565B;
wire g1918B;
wire g2340B;
wire g7684B;
wire g11519B;
wire g5935B;
wire g3800B;
wire g4736B;
wire g6941B;
wire g201B;
wire g2435B;
wire g4010B;
wire g1371B;
wire g2082B;
wire g4811B;
wire g5519B;
wire g49B;
wire g560B;
wire g6481B;
wire g6215B;
wire g10563B;
wire g10668B;
wire g70B;
wire g5013B;
wire g11221B;
wire g9508B;
wire g5212B;
wire g6529B;
wire g8709B;
wire g115B;
wire g2214B;
wire g5008B;
wire g3829B;
wire g9995B;
wire g10707B;
wire g3435B;
wire I7847B;
wire g5576B;
wire I13400B;
wire I5002B;
wire g10013B;
wire g10385B;
wire g9432B;
wire g3753B;
wire g4566B;
wire g254B;
wire I14326B;
wire g4722B;
wire g3348B;
wire g9696B;
wire g10408B;
wire I15968B;
wire g756B;
wire g818B;
wire g10937B;
wire g11060B;
wire g7242B;
wire g10336B;
wire I15855B;
wire g5229B;
wire g8940B;
wire g259B;
wire g10584B;
wire g10679B;
wire g4560B;
wire g10855B;
wire g369B;
wire g1968B;
wire I15503B;
wire g7996B;
wire g8110B;
wire g186B;
wire g2556B;
wire g3586B;
wire g10496B;
wire g3399B;
wire I7817B;
wire g158B;
wire g2222B;
wire g6907B;
wire g8226B;
wire I13373B;
wire g5405B;
wire I9880B;
wire g6155B;
wire g7246B;
wire g6638B;
wire g11647B;
wire g2744B;
wire g4094B;
wire g32B;
wire g3374B;
wire g4567B;
wire g8814B;
wire I14312B;
wire g10950B;
wire g9490B;
wire g11111B;
wire g4776B;
wire g5477B;
wire g6910B;
wire g10417B;
wire I15986B;
wire g713B;
wire g2237B;
wire g6488B;
wire g7712B;
wire g7897B;
wire g6828B;
wire g7638B;
wire g3015B;
wire g3121B;
wire I4917B;
wire g10800B;
wire g4300B;
wire g5420B;
wire g8019B;
wire I15956B;
wire g1840B;
wire g2557B;
wire g105B;
wire g9097B;
wire g6821B;
wire g3938B;
wire I5245B;
wire g253B;
wire g7682B;
wire g8267B;
wire g11478B;
wire g3698B;
wire g4379B;
wire g4144B;
wire g584B;
wire g131B;
wire g2254B;
wire g4289B;
wire g3992B;
wire g4777B;
wire I5424B;
wire g1776B;
wire g4585B;
wire g7934B;
wire g8089B;
wire g243B;
wire g2438B;
wire g6516B;
wire g8244B;
wire g4271B;
wire g4753B;
wire g8631B;
wire g4807B;
wire g10793B;
wire g7045B;
wire g5910B;
wire g9454B;
wire g686B;
wire g2212B;
wire I14299B;
wire g2563B;
wire g3141B;
wire g2478B;
wire g569B;
wire g35B;
wire g3215B;
wire g3710B;
wire I16252B;
wire g10726B;
wire g7516B;
wire g7920B;
wire g6824B;
wire g162B;
wire g2229B;
wire g9931B;
wire I15157B;
wire g11157B;
wire I15365B;
wire g79B;
wire I9279B;
wire g5361B;
wire g10558B;
wire g5248B;
wire g3880B;
wire g5557B;
wire g2172B;
wire g6759B;
wire g6502B;
wire g10797B;
wire g8241B;
wire I5044B;
wire g7685B;
wire g4471B;
wire g10780B;
wire g11625B;
wire g11372B;
wire g10007B;
wire I15287B;
wire g10771B;
wire I15290B;
wire g9720B;
wire g127B;
wire g2249B;
wire g5803B;
wire g11231B;
wire g11580B;
wire g5478B;
wire g11243B;
wire g4998B;
wire g10019B;
wire I5414B;
wire g4114B;
wire g11293B;
wire g2176B;
wire g4779B;
wire g5820B;
wire g8173B;
wire g3111B;
wire g3628B;
wire g4977B;
wire g6081B;
wire g255B;
wire g6533B;
wire I8503B;
wire g7460B;
wire g7910B;
wire g1984B;
wire g3688B;
wire g4285B;
wire g5867B;
wire g6354B;
wire g1690B;
wire g2031B;
wire g1857B;
wire I5510B;
wire g10405B;
wire g7932B;
wire g8085B;
wire g928B;
wire g7883B;
wire g10448B;
wire g5001B;
wire g8245B;
wire g3440B;
wire g4737B;
wire g8451B;
wire g8214B;
wire I13351B;
wire g3041B;
wire g10767B;
wire g10599B;
wire g10501B;
wire g3546B;
wire g8512B;
wire g2276B;
wire g6000B;
wire g6863B;
wire g10809B;
wire g10883B;
wire g5521B;
wire I14323B;
wire g11492B;
wire g932B;
wire g37B;
wire I6260B;
wire I9311B;
wire g4490B;
wire g8488B;
wire I5579B;
wire I9268B;
wire g4903B;
wire g10720B;
wire g10334B;
wire g10439B;
wire g6934B;
wire g5309B;
wire g5878B;
wire g4273B;
wire g7622B;
wire g6123B;
wire g7467B;
wire g774B;
wire g1990B;
wire g2248B;
wire g6838B;
wire g2045B;
wire g4905B;
wire g10798B;
wire g10785B;
wire g8187B;
wire I13436B;
wire g605B;
wire g2399B;
wire g7204B;
wire g6830B;
wire g6716B;
wire g8944B;
wire I5254B;
wire g5543B;
wire I5410B;
wire g5300B;
wire g8921B;
wire g8745B;
wire g8849B;
wire g6096B;
wire I7752B;
wire g6003B;
wire g3431B;
wire I7840B;
wire g10852B;
wire g6733B;
wire g7562B;
wire g6548B;
wire g1419B;
wire I9810B;
wire g5502B;
wire g260B;
wire g4679B;
wire g6823B;
wire g4890B;
wire g7981B;
wire g2579B;
wire g3776B;
wire g572B;
wire g3381B;
wire g10863B;
wire g971B;
wire g2008B;
wire g8039B;
wire g6526B;
wire g1900B;
wire g2336B;
wire g10664B;
wire g7189B;
wire g5278B;
wire g8923B;
wire g5173B;
wire g3521B;
wire I14306B;
wire g10712B;
wire I9296B;
wire g4264B;
wire g2178B;
wire g6755B;
wire g2791B;
wire I6962B;
wire g5226B;
wire g704B;
wire g2230B;
wire g4437B;
wire g11514B;
wire g7505B;
wire g38B;
wire g9507B;
wire g10411B;
wire I15974B;
wire g4506B;
wire g1834B;
wire g2550B;
wire g10348B;
wire g10400B;
wire I9282B;
wire I5584B;
wire g9324B;
wire g3664B;
wire g10001B;
wire g5526B;
wire g7697B;
wire g231B;
wire g2395B;
wire I5395B;
wire g4788B;
wire g4465B;
wire g8289B;
wire g6403B;
wire g8203B;
wire I15510B;
wire g5403B;
wire g6902B;
wire g6015B;
wire g11340B;
wire g6542B;
wire I5406B;
wire g3744B;
wire g581B;
wire I4883B;
wire g4537B;
wire g7688B;
wire g882B;
wire g2481B;
wire g6507B;
wire g10485B;
wire I4935B;
wire g10683B;
wire I9308B;
wire I5070B;
wire g5556B;
wire g8505B;
wire g8603B;
wire g11641B;
wire g3423B;
wire g4787B;
wire I9332B;
wire g10765B;
wire g6447B;
wire g4801B;
wire g11305B;
wire g3092B;
wire g6126B;
wire g4281B;
wire g5493B;
wire g5613B;
wire g639B;
wire g10414B;
wire g7986B;
wire g8255B;
wire g8000B;
wire g8081B;
wire g814B;
wire I9479B;
wire I4780B;
wire g2216B;
wire g10522B;
wire I5383B;
wire g8060B;
wire g7191B;
wire g8746B;
wire g8783B;
wire g10557B;
wire g5150B;
wire I5445B;
wire g4449B;
wire I4866B;
wire g6469B;
wire g7696B;
wire g10452B;
wire g4498B;
wire g8744B;
wire g8828B;
wire g2034B;
wire g2677B;
wire g5514B;
wire g6627B;
wire g4893B;
wire g10268B;
wire g10361B;
wire g3737B;
wire g9257B;
wire g9525B;
wire g5194B;
wire g668B;
wire g2198B;
wire g3418B;
wire I7771B;
wire g6901B;
wire g8043B;
wire g5263B;
wire g6929B;
wire g5857B;
wire g3523B;
wire g8049B;
wire g4529B;
wire g9699B;
wire g722B;
wire g2241B;
wire g6786B;
wire g7218B;
wire g7681B;
wire g6234B;
wire g5824B;
wire g7101B;
wire g10864B;
wire g7651B;
wire g7914B;
wire g986B;
wire I13427B;
wire g8816B;
wire I14319B;
wire I5430B;
wire g2175B;
wire g10862B;
wire I15980B;
wire g11077B;
wire I9259B;
wire g7683B;
wire I16717B;
wire I5388B;
wire I9326B;
wire g153B;
wire g2211B;
wire g3222B;
wire g3983B;
wire g4678B;
wire g3101B;
wire g3543B;
wire I5053B;
wire g9268B;
wire g5942B;
wire g10331B;
wire g10421B;
wire g10721B;
wire g8051B;
wire g2118B;
wire g10383B;
wire g6541B;
wire g936B;
wire g9088B;
wire g139B;
wire g2083B;
wire I6360B;
wire g10773B;
wire g8193B;
wire I4992B;
wire g6523B;
wire I16982B;
wire g8546B;
wire g8599B;
wire g794B;
wire g1828B;
wire g2061B;
wire g746B;
wire g2187B;
wire I9383B;
wire g5404B;
wire g11393B;
wire g5258B;
wire g1845B;
wire g2271B;
wire g1400B;
wire g2446B;
wire g8265B;
wire g2984B;
wire g11561B;
wire g11575B;
wire g822B;
wire g4765B;
wire g4334B;
wire g1936B;
wire g2345B;
wire g11233B;
wire g7950B;
wire g8106B;
wire g6586B;
wire g6908B;
wire g8768B;
wire g8885B;
wire g563B;
wire g33B;
wire g5808B;
wire I5418B;
wire g1361B;
wire g2016B;
wire g5271B;
wire g6333B;
wire g10515B;
wire g7692B;
wire I9273B;
wire g6045B;
wire g123B;
wire g731B;
wire g2251B;
wire g1988B;
wire g2047B;
wire g10927B;
wire g7590B;
wire g2275B;
wire g6468B;
wire g10782B;
wire g10886B;
wire g6672B;
wire g6840B;
wire g5230B;
wire g549B;
wire g8743B;
wire g8858B;
wire g3354B;
wire g4671B;
wire g5914B;
wire g7705B;
wire g7953B;
wire g8115B;
wire g10025B;
wire g1218B;
wire g2017B;
wire I5101B;
wire g6038B;
wire g1882B;
wire g2328B;
wire I5057B;
wire g1868B;
wire g2542B;
wire g4488B;
wire g1891B;
wire g2330B;
wire g3863B;
wire g6471B;
wire g11303B;
wire I9276B;
wire g7949B;
wire I5041B;
wire g782B;
wire g1992B;
wire I5441B;
wire g1110B;
wire g4365B;
wire g5266B;
wire g8234B;
wire I13364B;
wire g4158B;
wire g10663B;
wire g8920B;
wire g4283B;
wire I4859B;
wire g10788B;
wire g1397B;
wire g2456B;
wire g7512B;
wire g7919B;
wire g4484B;
wire I17413B;
wire I9346B;
wire g643B;
wire g1976B;
wire g7952B;
wire g865B;
wire I4820B;
wire I5435B;
wire g8815B;
wire I14315B;
wire g3008B;
wire g4467B;
wire g9713B;
wire g4290B;
wire g7527B;
wire g4770B;
wire g9474B;
wire g36B;
wire g5842B;
wire I9265B;
wire g7671B;
wire g8056B;
wire g8700B;
wire g4381B;
wire g5396B;
wire g1854B;
wire g7203B;
wire I6273B;
wire g10382B;
wire g10583B;
wire g10629B;
wire g8045B;
wire g7843B;
wire g2652B;
wire g754B;
wire g2057B;
wire g3539B;
wire g4263B;
wire g8269B;
wire I9349B;
wire I13323B;
wire g1386B;
wire g2549B;
wire g5261B;
wire g3104B;
wire g3419B;
wire g3425B;
wire I7829B;
wire g9802B;
wire g806B;
wire g6537B;
wire I13338B;
wire g5221B;
wire g3086B;
wire g2253B;
wire g4902B;
wire g6080B;
wire I9371B;
wire g5485B;
wire g6059B;
wire g4089B;
wire I5588B;
wire g7664B;
wire g7907B;
wire g4673B;
wire g8551B;
wire g5126B;
wire g10866B;
wire g10597B;
wire g11603B;
wire g6332B;
wire g4231B;
wire g9526B;
wire g207B;
wire g2570B;
wire g7473B;
wire g7915B;
wire I4783B;
wire g1991B;
wire g7677B;
wire g64B;
wire g11249B;
wire g636B;
wire g2506B;
wire g11348B;
wire g10779B;
wire g11488B;
wire g3491B;
wire g40B;
wire g3438B;
wire I7852B;
wire g757B;
wire g5354B;
wire g5295B;
wire g5918B;
wire g6894B;
wire g3513B;
wire g1713B;
wire I6240B;
wire g258B;
wire g591B;
wire g2374B;
wire g9424B;
wire g4076B;
wire g6534B;
wire g58B;
wire g3793B;
wire g6928B;
wire g7686B;
wire g3414B;
wire I7825B;
wire g8055B;
wire g11291B;
wire g237B;
wire g2420B;
wire g3209B;
wire g4739B;
wire g5509B;
wire g6833B;
wire g1958B;
wire g6918B;
wire g4608B;
wire I4948B;
wire g6915B;
wire g6911B;
wire I5060B;
wire g8812B;
wire I9237B;
wire g4553B;
wire g7441B;
wire g5996B;
wire g8047B;
wire g1786B;
wire g6653B;
wire g7438B;
wire g6832B;
wire I5047B;
wire g4771B;
wire g11481B;
wire g10857B;
wire g7947B;
wire g8100B;
wire g3681B;
wire g7918B;
wire I5427B;
wire g6478B;
wire g4117B;
wire g6897B;
wire g6042B;
wire I9717B;
wire g119B;
wire g11229B;
wire g1453B;
wire g2410B;
wire g10402B;
wire g4342B;
wire g4330B;
wire g8221B;
wire g1927B;
wire g2343B;
wire g11609B;
wire g10859B;
wire g6054B;
wire g6508B;
wire g6531B;
wire g8050B;
wire g8261B;
wire I9290B;
wire g11376B;
wire g580B;
wire I4876B;
wire g802B;
wire g8559B;
wire I9769B;
wire g2260B;
wire g10556B;
wire g148B;
wire g2202B;
wire g7032B;
wire g8390B;
wire g8548B;
wire g590B;
wire g2518B;
wire g4548B;
wire g4293B;
wire I16507B;
wire g5390B;
wire g4561B;
wire g8233B;
wire g1289B;
wire g8200B;
wire g4294B;
wire g76B;
wire g8767B;
wire g3071B;
wire g3723B;
wire I15962B;
wire g940B;
wire g7987B;
wire g8094B;
wire g1861B;
wire g2050B;
wire g1987B;
wire g4480B;
wire g11483B;
wire g1351B;
wire g10702B;
wire g5863B;
wire g2273B;
wire g5392B;
wire g9082B;
wire g5838B;
wire g8270B;
wire g10776B;
wire g2024B;
wire g2777B;
wire g6513B;
wire g9272B;
wire g10732B;
wire g1411B;
wire g10898B;
wire g869B;
wire g8052B;
wire g4325B;
wire g3368B;
wire g762B;
wire g4421B;
wire I8869B;
wire g5319B;
wire g8766B;
wire g10555B;
wire g586B;
wire g61B;
wire g6205B;
wire g778B;
wire g622B;
wire g8820B;
wire I9329B;
wire g11199B;
wire g9124B;
wire g6839B;
wire g6522B;
wire g10936B;
wire g7852B;
wire g7923B;
wire g11320B;
wire g6841B;
wire g10328B;
wire g10431B;
wire g8769B;
wire g6224B;
wire g2208B;
wire g11349B;
wire g4782B;
wire g6470B;
wire g11225B;
wire g5755B;
wire g4292B;
wire g1212B;
wire g6515B;
wire g3003B;
wire g3760B;
wire g9710B;
wire g5117B;
wire g3631B;
wire g5182B;
wire g11430B;
wire I9368B;
wire g10791B;
wire g5004B;
wire g1806B;
wire g7632B;
wire g11485B;
wire I5399B;
wire g6331B;
wire g1718B;
wire g2424B;
wire g5257B;
wire g8053B;
wire g4518B;
wire g7550B;
wire g219B;
wire g2077B;
wire g3103B;
wire g4764B;
wire g7913B;
wire g1989B;
wire g3068B;
wire g6109B;
wire I15500B;
wire g5763B;
wire g6480B;
wire g6795B;
wire g6449B;
wire g8194B;
wire g2257B;
wire g5201B;
wire g5269B;
wire g7497B;
wire g876B;
wire g2444B;
wire g1107B;
wire g8938B;
wire g7990B;
wire g8099B;
wire g4238B;
wire g8775B;
wire g4891B;
wire g8266B;
wire g11290B;
wire g6501B;
wire g10570B;
wire g10676B;
wire g6334B;
wire g786B;
wire g1993B;
wire g10719B;
wire g1104B;
wire g4727B;
wire g4274B;
wire g8765B;
wire g6916B;
wire g8811B;
wire I14303B;
wire g5174B;
wire I5525B;
wire I14330B;
wire g583B;
wire I4900B;
wire g11308B;
wire g3060B;
wire g5847B;
wire g10554B;
wire g10784B;
wire g2979B;
wire g599B;
wire g2382B;
wire g7680B;
wire g10396B;
wire g3784B;
wire g11425B;
wire I14295B;
wire g1346B;
wire I9293B;
wire I5815B;
wire g4002B;
wire g7062B;
wire g3479B;
wire g5548B;
wire g6131B;
wire g2449B;
wire g6820B;
wire g3390B;
wire g5627B;
wire g3501B;
wire g4340B;
wire I13385B;
wire g143B;
wire g2095B;
wire g1771B;
wire g257B;
wire g2297B;
wire g262B;
wire g6922B;
wire g1969B;
wire g6747B;
wire g11391B;
wire g8818B;
wire g8649B;
wire g9555B;
wire g6071B;
wire g1796B;
wire g7942B;
wire g8095B;
wire g6718B;
wire g611B;
wire g2364B;
wire g10858B;
wire g55B;
wire g1864B;
wire g2054B;
wire g2018B;
wire g2725B;
wire g627B;
wire g8926B;
wire g4239B;
wire g11602B;
wire g8041B;
wire g5503B;
wire g646B;
wire g1980B;
wire g981B;
wire g8164B;
wire g883B;
wire I6220B;
wire g582B;
wire I4891B;
wire g8922B;
wire g5536B;
wire g578B;
wire g5810B;
wire g7067B;
wire g8236B;
wire g11605B;
wire g8048B;
wire g6528B;
wire g1909B;
wire g2338B;
wire g34B;
wire g6524B;
wire g7446B;
wire g3056B;
wire g3475B;
wire g7258B;
wire g7219B;
wire g8046B;
wire g3706B;
wire g4822B;
wire g11482B;
wire g10381B;
wire g4477B;
wire g10333B;
wire g10437B;
wire g4456B;
wire g2310B;
wire g3039B;
wire g6923B;
wire g4255B;
wire g878B;
wire g790B;
wire g4732B;
wire g8937B;
wire g4752B;
wire g6538B;
wire g10339B;
wire g3524B;
wire g11306B;
wire g7183B;
wire g4778B;
wire g6165B;
wire g6895B;
wire g588B;
wire g11223B;
wire g6163B;
wire g6179B;
wire g9052B;
wire g9505B;
wire g9721B;
wire g654B;
wire g2268B;
wire g8776B;
wire g6827B;
wire g461B;
wire g4309B;
wire g9331B;
wire g7244B;
wire g7586B;
wire g7930B;
wire g5222B;
wire g11300B;
wire g10718B;
wire g213B;
wire g2070B;
wire g3906B;
wire g579B;
wire g5445B;
wire g11227B;
wire g6088B;
wire g658B;
wire g2331B;
wire g1365B;
wire g2406B;
wire g8206B;
wire I13332B;
wire g6679B;
wire g11636B;
wire g11239B;
wire g11219B;
wire g225B;
wire g2087B;
wire g2117B;
wire g2801B;
wire g3062B;
wire g3738B;
wire g9266B;
wire g9760B;
wire g11608B;
wire g8059B;
wire g8771B;
wire g2459B;
wire g6035B;
wire g1811B;
wire g7106B;
wire g471B;
wire g6198B;
wire g7992B;
wire g8105B;
wire g2169B;
wire g8973B;
wire g617B;
wire g2369B;
wire g6834B;
wire g197B;
wire g2407B;
wire g1962B;
wire g5148B;
wire I14642B;
wire g5836B;
wire g7134B;
wire I15514B;
wire g10795B;
wire g11083B;
wire g11276B;
wire g10770B;
wire g1810B;
wire g9271B;
wire g677B;
wire g2203B;
wire g587B;
wire I5497B;
wire I13421B;
wire g10494B;
wire g8773B;
wire g3462B;
wire I16220B;
wire g3662B;
wire g6740B;
wire g10484B;
wire g7143B;
wire g8939B;
wire g1703B;
wire g2028B;
wire g8772B;
wire g4336B;
wire g2067B;
wire g1814B;
wire g2564B;
wire g6093B;
wire g6500B;
wire g1407B;
wire g3705B;
wire g10500B;
wire g2794B;
wire g4065B;
wire g4243B;
wire g4934B;
wire g6485B;
wire g8777B;
wire g6244B;
wire g5304B;
wire g11640B;
wire g3814B;
wire g4784B;
wire g11487B;
wire g9110B;
wire g1822B;
wire g2571B;
wire g11380B;
wire g1950B;
wire g826B;
wire g9269B;
wire g7054B;
wire g1975B;
wire g7236B;
wire g2774B;
wire g3247B;
wire g3967B;
wire g11314B;
wire g585B;
wire g5276B;
wire g9150B;
wire g1389B;
wire g2396B;
wire g11298B;
wire g7202B;
wire g6819B;
wire g2987B;
wire g758B;
wire g11539B;
wire g1336B;
wire g108B;
wire g5317B;
wire g67B;
wire g10453B;
wire g6243B;
wire g6514B;
wire g8817B;
wire g8810B;
wire g1206B;
wire I6277B;
wire g1368B;
wire g2381B;
wire g9313B;
wire g10387B;
wire g6983B;
wire g8366B;
wire g8509B;
wire g7450B;
wire g7905B;
wire g4473B;
wire g6577B;
wire g1341B;
wire g1374B;
wire g2421B;
wire g3200B;
wire g4001B;
wire g8040B;
wire g5255B;
wire g6900B;
wire g8042B;
wire g11490B;
wire g11515B;
wire g8230B;
wire g6546B;
wire g3485B;
wire g1383B;
wire g2562B;
wire g6697B;
wire g8574B;
wire g5770B;
wire I11360B;
wire g8889B;
wire g10711B;
wire g9719B;
wire g11312B;
wire g5287B;
wire g11107B;
wire g1791B;
wire g6351B;
wire g9778B;
wire g6479B;
wire g3120B;
wire g3765B;
wire g5814B;
wire g5849B;
wire g1101B;
wire g575B;
wire g10559B;
wire g5219B;
wire g7240B;
wire I9352B;
wire g8819B;
wire g9256B;
wire g261B;
wire g6656B;
wire g976B;
wire g736B;
wire g1424B;
wire g1377B;
wire g2074B;
wire g6906B;
wire g10717B;
wire g4759B;
wire g5189B;
wire g8770B;
wire g6392B;
wire g6621B;
wire g11610B;
wire g4582B;
wire g6432B;
wire g7454B;
wire g7908B;
wire g8264B;
wire g11604B;
wire g9764B;
wire g2161B;
wire g3291B;
wire g7245B;
wire g2510B;
wire g256B;
wire g2439B;
wire g3207B;
wire g810B;
wire g11486B;
wire g12B;
wire g2126B;
wire g7581B;
wire g10799B;
wire I15507B;
wire I9221B;
wire g114B;
wire g1964B;
wire g10357B;
wire g6439B;
wire g8507B;
wire g8688B;
wire g7133B;
wire g8642B;
wire g8044B;
wire g8254B;
wire g11549B;
wire g1357B;
wire g2023B;
wire g7379B;
wire g11232B;
wire g11607B;
wire g6573B;
wire g3506B;
wire g3407B;
wire g770B;
wire g6193B;
wire g3108B;
wire g3408B;
wire g248B;
wire g2451B;
wire g7225B;
wire g8220B;
wire g7231B;
wire g4576B;
wire g3943B;
wire g4904B;
wire g8806B;
wire g11292B;
wire g6822B;
wire g7624B;
wire g3661B;
wire I15861B;
wire g73B;
wire g1801B;
wire g8327B;
wire g6912B;
wire g6898B;
wire g554B;
wire g8146B;
wire I5020B;
wire g5421B;
wire g1766B;
wire g7994B;
wire g8103B;
wire g1362B;
wire g2434B;
wire g3913B;
wire g6702B;
wire g4880B;
wire g8696B;
wire g868B;
wire g8813B;
wire I14309B;
wire g1945B;
wire g2347B;
wire g6924B;
wire g5308B;
wire g7574B;
wire g11310B;
wire g11294B;
wire g5852B;
wire g2970B;
wire g6026B;
wire g10369B;
wire g5286B;
wire g4554B;
wire g8024B;
wire g8945B;
wire g4804B;
wire g6525B;
wire g1380B;
wire g2060B;
wire g6019B;
wire g6617B;
wire g8210B;
wire g5083B;
wire g3585B;
wire g589B;
wire g7541B;
wire g4760B;
wire g26B;
wire g2479B;
wire g10860B;
wire g10502B;
wire g11579B;
wire g11639B;
wire g9814B;
wire g5030B;
wire g39B;
wire g6826B;
wire g2303B;
wire g9773B;
wire g52B;
wire g7626B;
wire g5200B;
wire g4457B;
wire g6829B;
wire g7211B;
wire g466B;
wire g456B;
wire g7660B;
wire g10722B;
wire g8887B;
wire g11484B;
wire g11286B;
wire g6002B;
wire g11606B;
wire g11217B;
wire g10454B;
wire g6757B;
wire g6216B;
wire g8941B;
wire g10856B;
wire g4892B;
wire g7903B;
wire g6930B;
wire g8250B;
wire g5250B;
wire g4525B;
wire g6049B;
wire g8943B;
wire g10861B;
wire g192B;
wire g2475B;
wire g8779B;
wire g766B;
wire g5484B;
wire g557B;
wire g11203B;
wire g3304B;
wire g6557B;
wire g4482B;
wire g1781B;
wire g5190B;
wire g6180B;
wire g5274B;
wire g8774B;
wire g10325B;
wire g10444B;
wire g566B;
wire g8260B;
wire g6099B;
wire g10401B;
wire g6831B;
wire g6068B;
wire g7137B;
wire g7917B;
wire g9473B;
wire g1965B;
wire g6545B;
wire g11547B;
wire g7257B;
wire g6909B;
wire g8384B;
wire g1872B;
wire g2503B;
wire g11392B;
wire g6506B;
wire g8883B;
wire g695B;
wire g2224B;
wire g6728B;
wire g10724B;
wire g4556B;
wire g3070B;
wire g2250B;
wire g11103B;
wire g9900B;
wire g845B;
wire g11095B;
wire g1645B;
wire g4973B;
wire g7389B;
wire g7465B;
wire g7888B;
wire g1642B;
wire g4969B;
wire g8224B;
wire g2892B;
wire g5686B;
wire g10308B;
wire g4123B;
wire g8120B;
wire g287B;
wire g6788B;
wire g4824B;
wire g5598B;
wire g278B;
wire g9694B;
wire g10495B;
wire g1684B;
wire g2945B;
wire g11190B;
wire g8639B;
wire g8789B;
wire g9728B;
wire g9563B;
wire g9852B;
wire g1053B;
wire g5625B;
wire g995B;
wire g4875B;
wire g1574B;
wire g9701B;
wire g7138B;
wire g10752B;
wire g11058B;
wire g11211B;
wire g435B;
wire g11024B;
wire g8307B;
wire g8547B;
wire g10669B;
wire g691B;
wire g7707B;
wire g3813B;
wire g4884B;
wire g4839B;
wire g1561B;
wire g9870B;
wire g6640B;
wire g9240B;
wire g9650B;
wire g5687B;
wire g7957B;
wire g3512B;
wire g7449B;
wire g1011B;
wire g4235B;
wire g345B;
wire g4343B;
wire g11296B;
wire g1B;
wire g9292B;
wire g9594B;
wire g1160B;
wire g9923B;
wire g9367B;
wire g9943B;
wire g1721B;
wire g5525B;
wire g440B;
wire g8876B;
wire g476B;
wire g10564B;
wire g10705B;
wire g9913B;
wire g9624B;
wire g9934B;
wire g6225B;
wire g1240B;
wire g6324B;
wire g10686B;
wire g1223B;
wire g6540B;
wire g8663B;
wire g1308B;
wire g11581B;
wire g6206B;
wire g452B;
wire g3989B;
wire g7260B;
wire g7730B;
wire g1235B;
wire g7504B;
wire g1887B;
wire g7185B;
wire I5689B;
wire I5690B;
wire g7881B;
wire g11070B;
wire g9736B;
wire g9859B;
wire g8877B;
wire g2274B;
wire g11590B;
wire g6199B;
wire g8932B;
wire g1730B;
wire g5545B;
wire g5180B;
wire g1615B;
wire g5591B;
wire g8412B;
wire g8556B;
wire g374B;
wire g11094B;
wire g5044B;
wire g5853B;
wire g6245B;
wire g4360B;
wire g8930B;
wire g5507B;
wire g3087B;
wire g11150B;
wire g8302B;
wire g8464B;
wire g272B;
wire g9692B;
wire g1428B;
wire g4996B;
wire g7131B;
wire g421B;
wire g11019B;
wire g9951B;
wire g9536B;
wire g9960B;
wire g11196B;
wire g11018B;
wire g10550B;
wire g10595B;
wire g10433B;
wire g10544B;
wire g10623B;
wire g4878B;
wire g4838B;
wire g5204B;
wire g8609B;
wire g8844B;
wire g6185B;
wire g6701B;
wire g10725B;
wire g5100B;
wire g1089B;
wire g4882B;
wire g8731B;
wire g1504B;
wire g5128B;
wire g1932B;
wire g6886B;
wire g8415B;
wire g8557B;
wire g8966B;
wire g8071B;
wire g11597B;
wire g9722B;
wire g9785B;
wire g9828B;
wire g1672B;
wire g2918B;
wire g9725B;
wire g9830B;
wire g8955B;
wire g4B;
wire g9592B;
wire g1618B;
wire g5123B;
wire g6078B;
wire g7059B;
wire g7459B;
wire g861B;
wire g11102B;
wire g709B;
wire g7718B;
wire g7535B;
wire g1577B;
wire g9703B;
wire g5528B;
wire g9911B;
wire g9932B;
wire g1636B;
wire g5530B;
wire g2760B;
wire g8629B;
wire g6187B;
wire g6887B;
wire g5605B;
wire g6228B;
wire g1275B;
wire g6322B;
wire I6337B;
wire I6338B;
wire g8967B;
wire g1458B;
wire g5010B;
wire g3275B;
wire g1678B;
wire g2895B;
wire g7721B;
wire g1549B;
wire g9866B;
wire g1534B;
wire g9716B;
wire g10744B;
wire g10808B;
wire g1231B;
wire g3047B;
wire g3685B;
wire g4492B;
wire g8614B;
wire g8822B;
wire g10560B;
wire g11456B;
wire g9724B;
wire g9848B;
wire g4714B;
wire g6550B;
wire g5172B;
wire g10642B;
wire g2531B;
wire g3284B;
wire g284B;
wire g302B;
wire g9855B;
wire g1630B;
wire g5618B;
wire g6891B;
wire g7940B;
wire g312B;
wire g11085B;
wire g396B;
wire g1432B;
wire g4968B;
wire g8646B;
wire g8837B;
wire g9125B;
wire g9644B;
wire g1546B;
wire g5804B;
wire g8300B;
wire g8462B;
wire I6330B;
wire g333B;
wire g11156B;
wire g293B;
wire g6342B;
wire g1552B;
wire g9867B;
wire g1537B;
wire g9717B;
wire g4871B;
wire g10435B;
wire g426B;
wire g7741B;
wire g1327B;
wire g9151B;
wire g9386B;
wire g8607B;
wire g8842B;
wire g8B;
wire g9599B;
wire g8974B;
wire g9274B;
wire g5518B;
wire g9111B;
wire g9614B;
wire g4122B;
wire g4610B;
wire g7217B;
wire g11557B;
wire g1675B;
wire g2911B;
wire g11210B;
wire g7466B;
wire g9918B;
wire g9939B;
wire g11279B;
wire g10513B;
wire g10440B;
wire I16145B;
wire g10518B;
wire g1129B;
wire g7055B;
wire g1095B;
wire g5264B;
wire g1265B;
wire g6329B;
wire g8176B;
wire g7510B;
wire g8005B;
wire g3281B;
wire g4099B;
wire g11601B;
wire g11187B;
wire g6746B;
wire g6221B;
wire g8630B;
wire g9622B;
wire g10923B;
wire g11143B;
wire g9886B;
wire g9676B;
wire g9904B;
wire g8733B;
wire g348B;
wire g6624B;
wire g530B;
wire g11169B;
wire g8073B;
wire g9706B;
wire g9512B;
wire g9841B;
wire g5592B;
wire g5882B;
wire g8645B;
wire g8796B;
wire g534B;
wire g11168B;
wire g1015B;
wire g4269B;
wire g727B;
wire g1047B;
wire g5611B;
wire g673B;
wire g8069B;
wire g1567B;
wire g9695B;
wire g10304B;
wire g8305B;
wire g8469B;
wire g1071B;
wire g4712B;
wire g5762B;
wire g6576B;
wire g10622B;
wire g5217B;
wire g11015B;
wire g5674B;
wire g9173B;
wire g9359B;
wire g8960B;
wire g9223B;
wire g11556B;
wire g1595B;
wire g9858B;
wire g5541B;
wire g363B;
wire g4534B;
wire g1499B;
wire g5897B;
wire g6177B;
wire g6699B;
wire g6855B;
wire g3098B;
wire g3804B;
wire g5680B;
wire g9642B;
wire g1528B;
wire g5744B;
wire g8399B;
wire g1762B;
wire g9030B;
wire g9447B;
wire g1849B;
wire g516B;
wire g11178B;
wire g8414B;
wire g8510B;
wire g1296B;
wire g6319B;
wire g11186B;
wire g1681B;
wire g2951B;
wire g6352B;
wire g9205B;
wire g9595B;
wire g4109B;
wire g4831B;
wire g1654B;
wire g5492B;
wire g8934B;
wire g10312B;
wire g6186B;
wire g9612B;
wire g1738B;
wire g9417B;
wire g9914B;
wire g9935B;
wire g10658B;
wire g10745B;
wire g956B;
wire g11216B;
wire g8971B;
wire g9328B;
wire g11587B;
wire g1245B;
wire g6325B;
wire g431B;
wire g7368B;
wire g552B;
wire g6083B;
wire g1227B;
wire g6544B;
wire g5476B;
wire g7743B;
wire g1083B;
wire g4869B;
wire g1598B;
wire g5722B;
wire g5813B;
wire g6790B;
wire g8408B;
wire g10761B;
wire g7734B;
wire g7926B;
wire g8136B;
wire g5569B;
wire g401B;
wire g9392B;
wire g9902B;
wire g8623B;
wire g1657B;
wire g5500B;
wire g2496B;
wire g3010B;
wire g5877B;
wire g6756B;
wire g8972B;
wire g336B;
wire g6622B;
wire g11612B;
wire g1311B;
wire g9366B;
wire g11230B;
wire g1284B;
wire g1215B;
wire g4364B;
wire g9649B;
wire g1543B;
wire g5795B;
wire g1524B;
wire g5737B;
wire g1753B;
wire g4054B;
wire g5823B;
wire g6345B;
wire g11275B;
wire g296B;
wire g9851B;
wire g5802B;
wire g6763B;
wire g416B;
wire g10511B;
wire g10509B;
wire g10507B;
wire I16142B;
wire g1571B;
wire g9698B;
wire g1032B;
wire g4725B;
wire g9954B;
wire g9964B;
wire g1663B;
wire g5523B;
wire g8402B;
wire g8550B;
wire g8611B;
wire g8845B;
wire g2081B;
wire g281B;
wire g6359B;
wire g1324B;
wire g11586B;
wire g5147B;
wire g11007B;
wire g5104B;
wire g4821B;
wire g5099B;
wire g5919B;
wire g1627B;
wire g5499B;
wire g3529B;
wire g4389B;
wire g3497B;
wire g6416B;
wire g1444B;
wire g4990B;
wire g9010B;
wire g9619B;
wire I6630B;
wire g6047B;
wire g953B;
wire g9652B;
wire g10505B;
wire g10469B;
wire g9711B;
wire g9519B;
wire g9843B;
wire g1074B;
wire g5273B;
wire g11465B;
wire g4348B;
wire g11237B;
wire g9731B;
wire g9834B;
wire g6654B;
wire g1041B;
wire g5444B;
wire g3714B;
wire g11285B;
wire g9598B;
wire g8097B;
wire g8726B;
wire g4816B;
wire g6880B;
wire g1157B;
wire g3287B;
wire g10759B;
wire g9917B;
wire g9938B;
wire g10652B;
wire g10758B;
wire g406B;
wire g9891B;
wire g9909B;
wire g6663B;
wire g7127B;
wire g11165B;
wire g1260B;
wire g6328B;
wire g8401B;
wire g5125B;
wire g11006B;
wire g1080B;
wire g4865B;
wire g1077B;
wire g4715B;
wire g2325B;
wire g4604B;
wire g5513B;
wire g965B;
wire g11222B;
wire g1145B;
wire g6554B;
wire g7732B;
wire g9586B;
wire g4401B;
wire g4104B;
wire g5178B;
wire g4584B;
wire g7472B;
wire g11253B;
wire g9860B;
wire g11600B;
wire g1586B;
wire g9645B;
wire g11236B;
wire g3106B;
wire g4162B;
wire g553B;
wire g6090B;
wire g269B;
wire g9691B;
wire g11316B;
wire g501B;
wire g11175B;
wire g664B;
wire g8068B;
wire g9607B;
wire g9952B;
wire g9962B;
wire g6348B;
wire g9659B;
wire g1318B;
wire g9358B;
wire I6316B;
wire I6317B;
wire g1711B;
wire g4486B;
wire g8995B;
wire g9587B;
wire g5632B;
wire g8965B;
wire g991B;
wire g4881B;
wire g11209B;
wire g8715B;
wire g8848B;
wire g3263B;
wire g4070B;
wire g6463B;
wire g1896B;
wire g7820B;
wire g448B;
wire g11021B;
wire g1044B;
wire g5917B;
wire g6619B;
wire g1300B;
wire g6318B;
wire g6872B;
wire g11201B;
wire g10489B;
wire g10514B;
wire g4006B;
wire g299B;
wire g9853B;
wire g11274B;
wire g8119B;
wire g1747B;
wire g9420B;
wire g5233B;
wire g7092B;
wire g6549B;
wire g11464B;
wire g4487B;
wire g1687B;
wire g2939B;
wire g6739B;
wire g7060B;
wire g1580B;
wire g5725B;
wire g11615B;
wire g2544B;
wire g11252B;
wire g5532B;
wire g3771B;
wire g11153B;
wire g9872B;
wire g9680B;
wire g9905B;
wire g7739B;
wire g6321B;
wire g8386B;
wire g8975B;
wire g2306B;
wire g6625B;
wire g7937B;
wire g8303B;
wire g8170B;
wire g5706B;
wire g2756B;
wire g8643B;
wire g8821B;
wire g5225B;
wire g10946B;
wire g4169B;
wire g5029B;
wire g11164B;
wire g4007B;
wire g1756B;
wire g4059B;
wire g1027B;
wire g4868B;
wire g5675B;
wire g4718B;
wire g10682B;
wire g6687B;
wire g682B;
wire g7704B;
wire g525B;
wire g1019B;
wire g4261B;
wire g3422B;
wire g5745B;
wire g8387B;
wire g7954B;
wire g11283B;
wire g8298B;
wire g8461B;
wire g10760B;
wire g11480B;
wire g6626B;
wire g6341B;
wire g10506B;
wire g16B;
wire g9648B;
wire g7453B;
wire g5995B;
wire g6645B;
wire g5707B;
wire g7548B;
wire g833B;
wire g11091B;
wire g496B;
wire g11174B;
wire g8403B;
wire g1250B;
wire g8605B;
wire g8841B;
wire g1914B;
wire g6879B;
wire g8763B;
wire g4502B;
wire g9702B;
wire g9839B;
wire g5841B;
wire g6358B;
wire g5575B;
wire g8107B;
wire g10240B;
wire g11192B;
wire g9618B;
wire g5539B;
wire g8416B;
wire g275B;
wire g9693B;
wire g11553B;
wire g7557B;
wire g1098B;
wire g5268B;
wire g9107B;
wire g10633B;
wire g7894B;
wire g8654B;
wire g9621B;
wire g5819B;
wire g6794B;
wire g3412B;
wire g7661B;
wire g2800B;
wire g3268B;
wire g9908B;
wire g3429B;
wire g351B;
wire g6628B;
wire g5470B;
wire g7526B;
wire g2204B;
wire g1482B;
wire g5025B;
wire g4921B;
wire g6204B;
wire g1750B;
wire g4048B;
wire g8935B;
wire g2525B;
wire g9593B;
wire g4827B;
wire g10701B;
wire g10733B;
wire g10777B;
wire g8130B;
wire g9955B;
wire g9965B;
wire g1710B;
wire g3684B;
wire g947B;
wire g11213B;
wire g1462B;
wire g5006B;
wire g9912B;
wire g9933B;
wire g8407B;
wire g8554B;
wire g9641B;
wire g6323B;
wire g10646B;
wire g10766B;
wire g6666B;
wire g4994B;
wire g5103B;
wire g3717B;
wire g11592B;
wire g1905B;
wire g6875B;
wire g9658B;
wire g6207B;
wire g6530B;
wire g8199B;
wire g7265B;
wire g9735B;
wire g9835B;
wire g6655B;
wire g3875B;
wire g7384B;
wire g7970B;
wire g1624B;
wire g5491B;
wire g8949B;
wire g11152B;
wire g9611B;
wire g2804B;
wire g6410B;
wire g10451B;
wire g4397B;
wire g5398B;
wire g7224B;
wire g5602B;
wire g6884B;
wire g8964B;
wire g11413B;
wire g1415B;
wire g4950B;
wire g5535B;
wire g6772B;
wire g7277B;
wire g8301B;
wire g8463B;
wire g2511B;
wire g10728B;
wire g6618B;
wire g6235B;
wire g6355B;
wire g3626B;
wire g4723B;
wire g8720B;
wire g6693B;
wire g11020B;
wire g1314B;
wire g11583B;
wire g8118B;
wire g8167B;
wire g7892B;
wire g8652B;
wire g5721B;
wire g10362B;
wire g10367B;
wire g9901B;
wire g290B;
wire g6792B;
wire g11282B;
wire g7945B;
wire g11302B;
wire g521B;
wire g3634B;
wire g11105B;
wire g8471B;
wire g8598B;
wire g7140B;
wire g9600B;
wire g1604B;
wire g9864B;
wire g11613B;
wire g5188B;
wire g7435B;
wire g7876B;
wire g1280B;
wire g4058B;
wire g5809B;
wire g6776B;
wire g630B;
wire g10301B;
wire g354B;
wire g4505B;
wire g17B;
wire g9623B;
wire g10739B;
wire g391B;
wire g11027B;
wire g10738B;
wire g8558B;
wire g8687B;
wire g6360B;
wire g1564B;
wire g9871B;
wire g5108B;
wire g11248B;
wire g4992B;
wire g11552B;
wire g944B;
wire g9651B;
wire g11204B;
wire g7824B;
wire g1133B;
wire g5115B;
wire g7102B;
wire g968B;
wire g9384B;
wire g2561B;
wire g9700B;
wire g9754B;
wire g9838B;
wire g10594B;
wire g10661B;
wire g11321B;
wire g8879B;
wire g7621B;
wire g8962B;
wire g2272B;
wire g10715B;
wire g8659B;
wire g950B;
wire g9643B;
wire g8957B;
wire g1669B;
wire g5538B;
wire g1744B;
wire g4000B;
wire g4126B;
wire g4088B;
wire g4400B;
wire I5886B;
wire I5887B;
wire g486B;
wire g6238B;
wire g10727B;
wire g8174B;
wire g305B;
wire g5067B;
wire g1512B;
wire g5418B;
wire g10297B;
wire g6353B;
wire g386B;
wire g11026B;
wire g11212B;
wire g4828B;
wire g6744B;
wire g1923B;
wire g10671B;
wire g2517B;
wire g4383B;
wire g4297B;
wire g5256B;
wire g4220B;
wire g8252B;
wire g8380B;
wire g7071B;
wire g9613B;
wire g8933B;
wire g5181B;
wire g7948B;
wire g324B;
wire g11149B;
wire g1601B;
wire g9862B;
wire g11387B;
wire g7955B;
wire g4161B;
wire g2321B;
wire g11148B;
wire g9712B;
wire g8931B;
wire g378B;
wire g11097B;
wire g3819B;
wire g2963B;
wire g11104B;
wire g1059B;
wire g6092B;
wire g4999B;
wire g4976B;
wire g632B;
wire g6858B;
wire g7409B;
wire g4103B;
wire I6309B;
wire g5944B;
wire g6580B;
wire g1056B;
wire g5631B;
wire g9414B;
wire g9660B;
wire g9926B;
wire g9946B;
wire I6331B;
wire g481B;
wire g9885B;
wire g9673B;
wire g9903B;
wire g10625B;
wire g6623B;
wire g11228B;
wire g11011B;
wire g1941B;
wire g6889B;
wire g7523B;
wire g7822B;
wire g8123B;
wire g11582B;
wire g4316B;
wire g3625B;
wire g10969B;
wire g5041B;
wire g9335B;
wire g9727B;
wire g9831B;
wire g9422B;
wire g4588B;
wire g8511B;
wire g8648B;
wire g8875B;
wire g5168B;
wire g7503B;
wire g7895B;
wire g8655B;
wire g1062B;
wire g4914B;
wire g9927B;
wire g9947B;
wire g1555B;
wire g5772B;
wire g1666B;
wire g5531B;
wire g5036B;
wire g10503B;
wire g7738B;
wire g8010B;
wire g8410B;
wire g5608B;
wire g6231B;
wire g10581B;
wire g10364B;
wire g10450B;
wire g2132B;
wire g2379B;
wire g9653B;
wire g1515B;
wire g10818B;
wire g8172B;
wire g10429B;
wire g5074B;
wire g1558B;
wire g9869B;
wire g10635B;
wire g10741B;
wire g8693B;
wire g5480B;
wire g3766B;
wire g4581B;
wire g2981B;
wire g8409B;
wire g8555B;
wire g9364B;
wire g506B;
wire g8994B;
wire g11299B;
wire g6592B;
wire g7958B;
wire g1474B;
wire g4995B;
wire g4079B;
wire g2264B;
wire g745B;
wire g2160B;
wire g3257B;
wire I6310B;
wire g1470B;
wire g5000B;
wire g3301B;
wire g1478B;
wire I5084B;
wire g1727B;
wire g9412B;
wire g1330B;
wire g9389B;
wire g10567B;
wire g10706B;
wire g10366B;
wire g10447B;
wire g10446B;
wire g10533B;
wire g5220B;
wire g10624B;
wire g10300B;
wire g5023B;
wire g4432B;
wire g4053B;
wire g7596B;
wire g1639B;
wire g5588B;
wire g6074B;
wire g9953B;
wire g9963B;
wire g3089B;
wire g3772B;
wire g5051B;
wire g8724B;
wire g4157B;
wire g1583B;
wire g9707B;
wire g8878B;
wire g10639B;
wire g10763B;
wire g6777B;
wire g8109B;
wire g7511B;
wire g7898B;
wire g11271B;
wire g11461B;
wire g5732B;
wire g315B;
wire g11145B;
wire g411B;
wire g11031B;
wire g1607B;
wire g9865B;
wire g1531B;
wire g9715B;
wire g9604B;
wire g8647B;
wire g8799B;
wire g11198B;
wire g6873B;
wire g6632B;
wire g6095B;
wire g9729B;
wire g9833B;
wire g1038B;
wire g6102B;
wire g7819B;
wire g11280B;
wire g7088B;
wire g9584B;
wire g9896B;
wire g8209B;
wire g6752B;
wire g11161B;
wire g8947B;
wire g5681B;
wire g7951B;
wire g9419B;
wire g1724B;
wire g5533B;
wire g8936B;
wire g178B;
wire g10670B;
wire g829B;
wire g11087B;
wire g4949B;
wire g5851B;
wire g6364B;
wire g7825B;
wire g1304B;
wire g10667B;
wire g7136B;
wire g339B;
wire g6532B;
wire g9385B;
wire g1436B;
wire g1440B;
wire g1448B;
wire g1137B;
wire g9897B;
wire g9425B;
wire g3383B;
wire g1035B;
wire g5601B;
wire g7943B;
wire g11171B;
wire I6631B;
wire g6064B;
wire g7230B;
wire g1648B;
wire g4952B;
wire g266B;
wire g6787B;
wire g8968B;
wire g10306B;
wire g11459B;
wire g538B;
wire g11458B;
wire g5739B;
wire g7496B;
wire g4986B;
wire g5187B;
wire g11010B;
wire g1741B;
wire g3999B;
wire g8175B;
wire g8722B;
wire g5590B;
wire g7471B;
wire g7891B;
wire g8651B;
wire g5479B;
wire g11599B;
wire g6684B;
wire g6745B;
wire g357B;
wire g6639B;
wire g3696B;
wire g4503B;
wire g6791B;
wire g8180B;
wire g1092B;
wire g4224B;
wire g5501B;
wire g8602B;
wire g8838B;
wire g10666B;
wire g309B;
wire g11158B;
wire g9602B;
wire g5704B;
wire g3879B;
wire g4617B;
wire g9868B;
wire g11295B;
wire g11144B;
wire g1540B;
wire g9718B;
wire g3434B;
wire g4987B;
wire g1270B;
wire g1065B;
wire g6098B;
wire g9582B;
wire g3533B;
wire g8104B;
wire g1733B;
wire g9415B;
wire g8377B;
wire g8499B;
wire g9664B;
wire g9413B;
wire g3584B;
wire g6162B;
wire g1508B;
wire g4991B;
wire g5846B;
wire g6362B;
wire g10685B;
wire g1153B;
wire g11023B;
wire g7598B;
wire g11224B;
wire g11571B;
wire g1520B;
wire g4959B;
wire g1633B;
wire g5626B;
wire g9920B;
wire g9940B;
wire g1086B;
wire g4876B;
wire g6730B;
wire g263B;
wire g9689B;
wire g10762B;
wire g1050B;
wire g6070B;
wire g9428B;
wire g1759B;
wire g9430B;
wire g8927B;
wire g7068B;
wire g7740B;
wire g8014B;
wire g11278B;
wire g5782B;
wire g4236B;
wire g11559B;
wire g9609B;
wire g11558B;
wire g6087B;
wire g10751B;
wire g10655B;
wire g10772B;
wire g8135B;
wire g11544B;
wire g5084B;
wire g8382B;
wire g10230B;
wire g7241B;
wire g3942B;
wire g10638B;
wire g4064B;
wire g1321B;
wire g9365B;
wire g9738B;
wire g9579B;
wire g9861B;
wire g11255B;
wire g11189B;
wire g10510B;
wire g2917B;
wire g11188B;
wire g9846B;
wire g1878B;
wire g7818B;
wire g11460B;
wire g11030B;
wire g841B;
wire g11093B;
wire g7478B;
wire g7893B;
wire g8653B;
wire g10442B;
wire g6535B;
wire g8102B;
wire g1490B;
wire g1494B;
wire I5085B;
wire g3912B;
wire g7186B;
wire g4489B;
wire g9662B;
wire g9418B;
wire g959B;
wire g11218B;
wire g1121B;
wire g10643B;
wire g10746B;
wire g7125B;
wire g7821B;
wire g6246B;
wire g8963B;
wire g7533B;
wire g10237B;
wire g7939B;
wire g8638B;
wire g8786B;
wire g10684B;
wire g11455B;
wire g8364B;
wire g2990B;
wire g9847B;
wire g7584B;
wire g5617B;
wire g5981B;
wire g5789B;
wire g4009B;
wire g11277B;
wire g6472B;
wire g6940B;
wire g6760B;
wire g7061B;
wire g11595B;
wire g5771B;
wire g8405B;
wire g8553B;
wire g4836B;
wire g5547B;
wire g4967B;
wire g342B;
wire g6671B;
wire g7200B;
wire g382B;
wire g7046B;
wire g999B;
wire g4229B;
wire g8389B;
wire g6430B;
wire g4993B;
wire g6247B;
wire g11170B;
wire g7145B;
wire g5738B;
wire g3998B;
wire g6741B;
wire g11167B;
wire g11194B;
wire g1333B;
wire g11589B;
wire g4431B;
wire g7536B;
wire g9585B;
wire g2957B;
wire g11588B;
wire g5690B;
wire g6883B;
wire g1068B;
wire g4837B;
wire g8641B;
wire g8791B;
wire g6217B;
wire g444B;
wire g11022B;
wire g4168B;
wire g5915B;
wire g511B;
wire g5110B;
wire g11254B;
wire g7567B;
wire g3273B;
wire g4392B;
wire g1592B;
wire g9856B;
wire g9411B;
wire g5002B;
wire g857B;
wire g11101B;
wire g11177B;
wire g11560B;
wire g8098B;
wire g3970B;
wire g4941B;
wire g366B;
wire g6662B;
wire g7935B;
wire g6067B;
wire g9740B;
wire g9863B;
wire g174B;
wire g170B;
wire g6758B;
wire g6994B;
wire g1589B;
wire g1007B;
wire g4252B;
wire g542B;
wire g11166B;
wire g7130B;
wire g5179B;
wire g11009B;
wire g7542B;
wire g5171B;
wire g11008B;
wire g1209B;
wire g3516B;
wire g7573B;
wire g3987B;
wire g491B;
wire g11555B;
wire g9734B;
wire g9569B;
wire g9857B;
wire g8728B;
wire g8730B;
wire g8185B;
wire g1610B;
wire g8385B;
wire g7902B;
wire g4073B;
wire g8070B;
wire g5731B;
wire g11238B;
wire g1125B;
wire g8308B;
wire g8470B;
wire g5489B;
wire g3991B;
wire g166B;
wire g7823B;
wire g4069B;
wire g1317B;
wire g11176B;
wire g837B;
wire g11092B;
wire g330B;
wire g11154B;
wire g7B;
wire g9608B;
wire g11637B;
wire g2091B;
wire g8406B;
wire g5254B;
wire g8612B;
wire g9588B;
wire g8742B;
wire g8801B;
wire g7063B;
wire g10303B;
wire g1486B;
wire g5009B;
wire g9665B;
wire g8748B;
wire g11215B;
wire g10750B;
wire g3818B;
wire g5769B;
wire g6673B;
wire g1255B;
wire g7720B;
wire g4609B;
wire g7547B;
wire g7971B;
wire g11288B;
wire g7599B;
wire g6058B;
wire g4106B;
wire g6743B;
wire g6890B;
wire g7269B;
wire g7549B;
wire g8169B;
wire g11304B;
wire g9924B;
wire g9944B;
wire g7592B;
wire g8718B;
wire g8616B;
wire g9316B;
wire g7625B;
wire g8644B;
wire g8793B;
wire g2940B;
wire g11624B;
wire g2947B;
wire g10949B;
wire g3563B;
wire g2223B;
wire g10948B;
wire g7846B;
wire g8246B;
wire g5788B;
wire g4008B;
wire g9596B;
wire g5249B;
wire g11585B;
wire g4972B;
wire g11554B;
wire g7096B;
wire g10673B;
wire g2493B;
wire g4806B;
wire g9915B;
wire g9936B;
wire g1660B;
wire g2910B;
wire g9317B;
wire g10853B;
wire g10933B;
wire g8177B;
wire g8388B;
wire g1117B;
wire g7141B;
wire g10508B;
wire g4230B;
wire g10634B;
wire g9192B;
wire g9601B;
wire g6326B;
wire g700B;
wire g7710B;
wire g7375B;
wire g8028B;
wire g5640B;
wire g5031B;
wire g4550B;
wire g7879B;
wire g7962B;
wire g9597B;
wire g631B;
wire g5005B;
wire g6423B;
wire g8108B;
wire g3322B;
wire g5911B;
wire g9916B;
wire g9937B;
wire g9704B;
wire g9747B;
wire g9840B;
wire g10723B;
wire g8217B;
wire g5209B;
wire g11013B;
wire g9390B;
wire g11214B;
wire g6327B;
wire g1149B;
wire g5796B;
wire g5473B;
wire g5038B;
wire g6346B;
wire g6633B;
wire g5119B;
wire g11005B;
wire g8365B;
wire g7558B;
wire g4481B;
wire g4097B;
wire g7588B;
wire g4497B;
wire g9922B;
wire g9942B;
wire g6696B;
wire g5118B;
wire g1850B;
wire g10665B;
wire g10731B;
wire g8552B;
wire g8827B;
wire g5540B;
wire g1403B;
wire g4960B;
wire g8615B;
wire g8846B;
wire g5983B;
wire g182B;
wire g6240B;
wire g7931B;
wire g853B;
wire g11100B;
wire g11235B;
wire g5199B;
wire g6316B;
wire g7515B;
wire g5781B;
wire g7742B;
wire g8018B;
wire g2950B;
wire g5510B;
wire g6347B;
wire g962B;
wire g9357B;
wire g11407B;
wire g10743B;
wire g5259B;
wire g5694B;
wire g10769B;
wire g11584B;
wire g4932B;
wire g10649B;
wire g10768B;
wire g4068B;
wire g6317B;
wire g4276B;
wire g5215B;
wire g6775B;
wire g10662B;
wire g8101B;
wire g3204B;
wire g5318B;
wire g5825B;
wire g7457B;
wire g7884B;
wire g1292B;
wire g3974B;
wire g9929B;
wire g9949B;
wire g10778B;
wire g7524B;
wire g6079B;
wire g7235B;
wire g9603B;
wire g9726B;
wire g9850B;
wire g7988B;
wire g5228B;
wire g5587B;
wire g5934B;
wire g8168B;
wire g9583B;
wire g10672B;
wire g8627B;
wire g635B;
wire g8309B;
wire g10449B;
wire g11273B;
wire g8734B;
wire g5913B;
wire g4572B;
wire g6363B;
wire g11463B;
wire g718B;
wire g8074B;
wire g1166B;
wire g8383B;
wire g8474B;
wire g11234B;
wire g4483B;
wire g11491B;
wire g5097B;
wire g5726B;
wire g5497B;
wire g7933B;
wire g9B;
wire g9617B;
wire g9873B;
wire g9906B;
wire g5196B;
wire g11012B;
wire g7050B;
wire g10849B;
wire g10971B;
wire g8400B;
wire g1169B;
wire g4345B;
wire g9925B;
wire g9945B;
wire g5028B;
wire g7271B;
wire g9709B;
wire g1003B;
wire g4223B;
wire g10497B;
wire g10716B;
wire g11247B;
wire g6661B;
wire g11173B;
wire g6075B;
wire g7367B;
wire g8023B;
wire g9888B;
wire g9907B;
wire g10582B;
wire g5746B;
wire g9950B;
wire g9959B;
wire g7674B;
wire g9690B;
wire g5703B;
wire g360B;
wire g4522B;
wire g4115B;
wire g7075B;
wire g10627B;
wire g4047B;
wire g2944B;
wire g6646B;
wire g7132B;
wire g11029B;
wire g7572B;
wire g8127B;
wire g7209B;
wire g11028B;
wire g10742B;
wire g8880B;
wire g10681B;
wire g9663B;
wire g5349B;
wire g8732B;
wire g3807B;
wire g3860B;
wire g5848B;
wire g8411B;
wire g8508B;
wire g8072B;
wire g5699B;
wire g11240B;
wire g6105B;
wire g6616B;
wire g10690B;
wire g7582B;
wire g9590B;
wire g4128B;
wire g6404B;
wire g6647B;
wire g10504B;
wire g9657B;
wire g4542B;
wire g1163B;
wire g5524B;
wire g9899B;
wire g7736B;
wire g10626B;
wire g6320B;
wire g7623B;
wire g10299B;
wire g7889B;
wire g10298B;
wire g8413B;
wire g3979B;
wire g1848B;
wire g5211B;
wire g4512B;
wire g7722B;
wire g9714B;
wire g9522B;
wire g9844B;
wire g1141B;
wire g5993B;
wire g5026B;
wire g8705B;
wire g10737B;
wire g10232B;
wire g6771B;
wire g5170B;
wire g8117B;
wire g9956B;
wire g9966B;
wire g5280B;
wire g7139B;
wire g11099B;
wire g6892B;
wire g9705B;
wire g10512B;
wire g849B;
wire g11098B;
wire g8628B;
wire g5544B;
wire g11272B;
wire g1621B;
wire g5483B;
wire g9928B;
wire g9948B;
wire g4063B;
wire g11462B;
wire g6738B;
wire g7593B;
wire g11032B;
wire g10445B;
wire g8882B;
wire g10316B;
wire g5756B;
wire g1023B;
wire g4720B;
wire g9409B;
wire g8929B;
wire g6876B;
wire g4989B;
wire g9737B;
wire g9836B;
wire g6061B;
wire g8268B;
wire g6465B;
wire g1466B;
wire g5003B;
wire g9957B;
wire g9967B;
wire g5145B;
wire g4971B;
wire g10753B;
wire g5695B;
wire g7613B;
wire g10736B;
wire g11220B;
wire g7444B;
wire g4670B;
wire g4253B;
wire g7960B;
wire g8163B;
wire g10764B;
wire g5757B;
wire g7385B;
wire g8032B;
wire g2988B;
wire g11591B;
wire g7583B;
wire g321B;
wire g11147B;
wire g5522B;
wire g1394B;
wire g9697B;
wire g9751B;
wire g9837B;
wire g9620B;
wire g327B;
wire g11151B;
wire g11172B;
wire g7885B;
wire g5595B;
wire g5537B;
wire g9708B;
wire g9516B;
wire g9842B;
wire g4141B;
wire g4341B;
wire g7679B;
wire g7378B;
wire g5612B;
wire g7135B;
wire g10970B;
wire g11025B;
wire g9730B;
wire g9854B;
wire g7182B;
wire g9921B;
wire g9941B;
wire g6194B;
wire g1651B;
wire g4962B;
wire g4358B;
wire g4803B;
wire g8549B;
wire g8683B;
wire g1113B;
wire g5224B;
wire g8778B;
wire g11281B;
wire g318B;
wire g11146B;
wire g2948B;
wire g3904B;
wire g8075B;
wire g9723B;
wire g9829B;
wire g7184B;
wire g11246B;
wire g5837B;
wire g6350B;
wire g2555B;
wire g5902B;
wire g1765B;
wire g6438B;
wire g5512B;
wire g5090B;
wire g7719B;
wire g3695B;
wire g7587B;
wire g9610B;
wire g3536B;
wire g8881B;
wire g4559B;
wire g10549B;
wire g10561B;
wire g5698B;
wire g11226B;
wire g10295B;
wire g5260B;
wire g10680B;
wire g1853B;
wire g11538B;
wire g11551B;
wire g9849B;
wire g5279B;
wire g8404B;
wire g5720B;
wire g11318B;
wire g11297B;
wire g9898B;
wire g9510B;
wire g7297B;
wire g7963B;
wire g9759B;
wire g9803B;
wire g11338B;
wire g8435B;
wire g6124B;
wire I5600B;
wire g11257B;
wire g11256B;
wire g3107B;
wire g2167B;
wire I14866B;
wire g4997B;
wire g10291B;
wire g6122B;
wire g9509B;
wire g5227B;
wire I15054B;
wire g11269B;
wire g5555B;
wire g11268B;
wire g11335B;
wire g8249B;
wire g9882B;
wire I15210B;
wire g2102B;
wire g2099B;
wire g2096B;
wire g2088B;
wire I5805B;
wire g11443B;
wire g8431B;
wire g8286B;
wire g7290B;
wire g8287B;
wire g7301B;
wire g8259B;
wire g11334B;
wire g10805B;
wire I15214B;
wire I15215B;
wire g11265B;
wire g8322B;
wire g8433B;
wire g8248B;
wire g8154B;
wire g2405B;
wire g2389B;
wire g2380B;
wire g2372B;
wire I6351B;
wire I16427B;
wire g7303B;
wire g2862B;
wire g2515B;
wire g4052B;
wire I14858B;
wire g11264B;
wire I15209B;
wire g1570B;
wire g2528B;
wire g2522B;
wire g9515B;
wire g7294B;
wire g3118B;
wire g2180B;
wire I5571B;
wire I5599B;
wire g2514B;
wire g11327B;
wire I5629B;
wire I5363B;
wire g2315B;
wire g8159B;
wire g11326B;
wire I16148B;
wire I16149B;
wire g10521B;
wire g7292B;
wire g8417B;
wire I14855B;
wire g9878B;
wire I15205B;
wire I15051B;
wire g8823B;
wire g8148B;
wire g2863B;
wire g2516B;
wire g7299B;
wire g9511B;
wire g9654B;
wire I15224B;
wire I15225B;
wire g8253B;
wire I15171B;
wire I15172B;
wire I15204B;
wire g10472B;
wire g10470B;
wire g10468B;
wire g10467B;
wire g10386B;
wire g10384B;
wire g10476B;
wire g10474B;
wire g8158B;
wire g11331B;
wire g7295B;
wire g8284B;
wire g1393B;
wire I5357B;
wire g9758B;
wire I5626B;
wire g7298B;
wire g8282B;
wire I15057B;
wire I15219B;
wire I15220B;
wire I14862B;
wire g2521B;
wire g9591B;
wire g9757B;
wire g11261B;
wire g9815B;
wire I14835B;
wire g126B;
wire g10479B;
wire g10478B;
wire g10477B;
wire g10475B;
wire I16161B;
wire g2353B;
wire I5804B;
wire g7291B;
wire I15199B;
wire g11330B;
wire g8153B;
wire g9881B;
wire g11259B;
wire g11258B;
wire g9426B;
wire g9423B;
wire g11337B;
wire g8262B;
wire g8285B;
wire I5570B;
wire g2499B;
wire g11336B;
wire g7293B;
wire g9388B;
wire g11260B;
wire g10807B;
wire g8288B;
wire g10394B;
wire g10392B;
wire g10482B;
wire g10481B;
wire I16160B;
wire g9589B;
wire g11270B;
wire g11267B;
wire g1959B;
wire g9667B;
wire I14827B;
wire g9391B;
wire I5358B;
wire g2309B;
wire g11266B;
wire g8429B;
wire g8281B;
wire g9876B;
wire I15177B;
wire g5186B;
wire I6350B;
wire g1527B;
wire g8162B;
wire I14779B;
wire I5351B;
wire I5352B;
wire g2305B;
wire I15176B;
wire g9879B;
wire g8283B;
wire g11333B;
wire g10562B;
wire g9606B;
wire I14822B;
wire g9880B;
wire I15200B;
wire g8428B;
wire g8430B;
wire g8247B;
wire I5576B;
wire g4476B;
wire I5649B;
wire g2538B;
wire g11329B;
wire g11328B;
wire g9605B;
wire g9363B;
wire g7300B;
wire I14831B;
wire g8263B;
wire g11263B;
wire g5780B;
wire g11332B;
wire I15048B;
wire g9647B;
wire I14602B;
wire I15033B;
wire g2445B;
wire g2437B;
wire g2433B;
wire g2419B;
wire g11325B;
wire I5366B;
wire g9506B;
wire g8161B;
wire g2316B;
wire g4675B;
wire g8434B;
wire g11262B;
wire g9387B;
wire I15045B;
wire g11324B;
wire g2501B;
wire g9877B;
wire g10529B;
wire g8432B;
wire g9874B;
wire g8157B;
wire g6899B;
wire g9646B;
wire g7302B;
wire g2111B;
wire g2109B;
wire g2106B;
wire g2104B;
wire g7296B;
wire I5612B;
wire I5613B;
wire I5591B;
wire I5593B;
wire g8839B;
wire g8970B;
wire I10519B;
wire I11278B;
wire I11279B;
wire g3978B;
wire I5263B;
wire I5264B;
wire g4278B;
wire I8640B;
wire g2943B;
wire I6760B;
wire I6761B;
wire g11418B;
wire g11416B;
wire I17400B;
wire I5449B;
wire I5450B;
wire I16058B;
wire I16060B;
wire g2938B;
wire I6746B;
wire I11973B;
wire I11975B;
wire I12136B;
wire I11935B;
wire I11937B;
wire I6167B;
wire I6168B;
wire g2959B;
wire g2120B;
wire g2115B;
wire I5878B;
wire I5619B;
wire I5620B;
wire g5552B;
wire I6467B;
wire I6468B;
wire g4672B;
wire I8795B;
wire I8796B;
wire I15891B;
wire I15892B;
wire I5611B;
wire g8738B;
wire I6714B;
wire I6716B;
wire g3460B;
wire I7683B;
wire I7685B;
wire I12106B;
wire I12108B;
wire I6747B;
wire I5230B;
wire I5231B;
wire g2236B;
wire I12075B;
wire I12076B;
wire I15870B;
wire I16065B;
wire I16067B;
wire I7562B;
wire I13529B;
wire I13531B;
wire I8797B;
wire I17584B;
wire I11936B;
wire I15256B;
wire I15257B;
wire I13505B;
wire I13506B;
wire g8502B;
wire g8501B;
wire g8824B;
wire I6186B;
wire I17504B;
wire I17505B;
wire g11496B;
wire I15999B;
wire I16001B;
wire g2215B;
wire I6124B;
wire I6125B;
wire I11907B;
wire I11909B;
wire I12038B;
wire I12040B;
wire I13907B;
wire I13909B;
wire I6771B;
wire I6772B;
wire I11908B;
wire I16008B;
wire I16009B;
wire I13908B;
wire I7034B;
wire I7035B;
wire I8650B;
wire I9947B;
wire I9948B;
wire g10428B;
wire I16066B;
wire I6144B;
wire I6145B;
wire I11241B;
wire I11242B;
wire I15993B;
wire I15994B;
wire I6187B;
wire g6027B;
wire I5500B;
wire I11974B;
wire I12060B;
wire I12062B;
wire I8771B;
wire I8772B;
wire I5184B;
wire I13293B;
wire I6199B;
wire I6200B;
wire I13265B;
wire I5023B;
wire I5024B;
wire I7863B;
wire I13991B;
wire I13992B;
wire I13660B;
wire I13661B;
wire I6143B;
wire I13990B;
wire I11508B;
wire I11510B;
wire g5034B;
wire I5229B;
wire I12045B;
wire I12047B;
wire I10769B;
wire I10771B;
wire I16045B;
wire I16046B;
wire I12061B;
wire I5104B;
wire I13530B;
wire I6447B;
wire I4954B;
wire I4956B;
wire g3530B;
wire I8479B;
wire I8481B;
wire I8739B;
wire I8740B;
wire I6879B;
wire I6880B;
wire I15430B;
wire I15431B;
wire I12019B;
wire I12020B;
wire I16331B;
wire I16332B;
wire I16467B;
wire I16469B;
wire I5013B;
wire I5014B;
wire I13521B;
wire I13523B;
wire I16037B;
wire I16039B;
wire I16468B;
wire I12046B;
wire I16038B;
wire g4374B;
wire I8676B;
wire I12113B;
wire g4616B;
wire I8761B;
wire I15992B;
wire I5034B;
wire I5036B;
wire g8843B;
wire I14263B;
wire I13249B;
wire I13250B;
wire I5135B;
wire I5485B;
wire I5486B;
wire I7033B;
wire I15441B;
wire I15443B;
wire I6166B;
wire g4267B;
wire I8624B;
wire I16015B;
wire I8677B;
wire g4234B;
wire I8575B;
wire I8576B;
wire g9204B;
wire I14612B;
wire I14613B;
wire g4601B;
wire I8715B;
wire I8716B;
wire I6715B;
wire I13514B;
wire I13515B;
wire I12002B;
wire I12003B;
wire I5127B;
wire I5128B;
wire g2177B;
wire I8577B;
wire g11414B;
wire I17393B;
wire I17395B;
wire I11280B;
wire I5265B;
wire I6988B;
wire I6989B;
wire I13272B;
wire I13274B;
wire I10507B;
wire I5164B;
wire I14443B;
wire I14444B;
wire I9557B;
wire I9559B;
wire I5592B;
wire I13077B;
wire I13078B;
wire I8717B;
wire I5295B;
wire I5296B;
wire I8625B;
wire I8626B;
wire I4911B;
wire I4912B;
wire I16000B;
wire I5371B;
wire I5185B;
wire I5186B;
wire I5675B;
wire g4218B;
wire I8543B;
wire I8544B;
wire I10520B;
wire I10521B;
wire I5297B;
wire I13537B;
wire I13283B;
wire g4749B;
wire I11980B;
wire I11982B;
wire g4873B;
wire I8513B;
wire I8514B;
wire I13089B;
wire I13091B;
wire I6126B;
wire g10302B;
wire I15906B;
wire I15908B;
wire I8763B;
wire g8506B;
wire g8825B;
wire I16007B;
wire g2107B;
wire g2105B;
wire I5865B;
wire I5604B;
wire I5517B;
wire I5518B;
wire I6109B;
wire I6111B;
wire I4929B;
wire I4930B;
wire I13522B;
wire I10770B;
wire I5538B;
wire I5539B;
wire g11415B;
wire I17394B;
wire I13552B;
wire I13553B;
wire I8642B;
wire I17296B;
wire I17297B;
wire I14278B;
wire I14279B;
wire I4910B;
wire I6792B;
wire I6794B;
wire I5484B;
wire I15442B;
wire I10931B;
wire I10932B;
wire I8779B;
wire I8780B;
wire g2354B;
wire g10043B;
wire g10153B;
wire I15615B;
wire I17281B;
wire I5468B;
wire I5470B;
wire I11509B;
wire I5025B;
wire I14270B;
wire I14272B;
wire I6208B;
wire I6209B;
wire I17288B;
wire I17290B;
wire I7563B;
wire I7564B;
wire I5005B;
wire I5006B;
wire I12126B;
wire I12128B;
wire I5105B;
wire I6322B;
wire I6323B;
wire I12093B;
wire I12094B;
wire g2776B;
wire I6664B;
wire I6666B;
wire I6762B;
wire g3623B;
wire I5373B;
wire I8527B;
wire I8529B;
wire I5282B;
wire I5283B;
wire I7223B;
wire I7224B;
wire I5007B;
wire I5459B;
wire I17295B;
wire I5015B;
wire I14264B;
wire I14265B;
wire I16072B;
wire I16073B;
wire g3205B;
wire I8652B;
wire I9558B;
wire I5202B;
wire I5203B;
wire I6806B;
wire I6807B;
wire I6469B;
wire I12143B;
wire I12145B;
wire I12127B;
wire I13300B;
wire I13302B;
wire I5502B;
wire I9574B;
wire I6448B;
wire I6449B;
wire I8669B;
wire I8670B;
wire I15451B;
wire I15453B;
wire I7875B;
wire I7876B;
wire I14202B;
wire I14203B;
wire g10149B;
wire g10144B;
wire I15607B;
wire I5324B;
wire I5325B;
wire I8738B;
wire g10434B;
wire g5859B;
wire I8604B;
wire I8606B;
wire I12085B;
wire I12087B;
wire I13248B;
wire I4979B;
wire I4980B;
wire I12067B;
wire I12069B;
wire g8942B;
wire I12068B;
wire I17503B;
wire I7877B;
wire I5165B;
wire I6287B;
wire I6289B;
wire I6777B;
wire I8562B;
wire I8563B;
wire I15890B;
wire g8006B;
wire I13090B;
wire I17460B;
wire I17461B;
wire g11474B;
wire I13513B;
wire I4986B;
wire I4987B;
wire I5204B;
wire I13504B;
wire I6207B;
wire I12086B;
wire I8545B;
wire I8178B;
wire I8180B;
wire I8589B;
wire I8591B;
wire I10930B;
wire I17402B;
wire I13294B;
wire I13295B;
wire I12144B;
wire g8757B;
wire g2961B;
wire I14209B;
wire I14211B;
wire I8515B;
wire I5316B;
wire I5317B;
wire I9946B;
wire g4613B;
wire I8750B;
wire I5605B;
wire I14204B;
wire I16051B;
wire g10360B;
wire g6037B;
wire I13858B;
wire I13859B;
wire I15872B;
wire g4879B;
wire I8528B;
wire I13901B;
wire I13902B;
wire g8542B;
wire I6836B;
wire I6838B;
wire I17305B;
wire I17307B;
wire g4538B;
wire I15452B;
wire I13857B;
wire I13765B;
wire I8671B;
wire I16044B;
wire g10363B;
wire g5360B;
wire I5106B;
wire g4677B;
wire I8803B;
wire I8804B;
wire I16016B;
wire I16017B;
wire I17485B;
wire I17487B;
wire I4995B;
wire I12092B;
wire I8678B;
wire I5126B;
wire I5372B;
wire I17306B;
wire I11995B;
wire I7225B;
wire I11261B;
wire g8545B;
wire I6110B;
wire I4941B;
wire I4942B;
wire I15899B;
wire I15900B;
wire g5527B;
wire g5350B;
wire I16079B;
wire I16081B;
wire I8641B;
wire I6176B;
wire I6178B;
wire I12074B;
wire I5451B;
wire I7322B;
wire I7323B;
wire I6288B;
wire I8179B;
wire I6805B;
wire I17486B;
wire I4928B;
wire I16330B;
wire I9575B;
wire I13886B;
wire I13887B;
wire I8787B;
wire I8788B;
wire I5315B;
wire g10285B;
wire I13867B;
wire I13869B;
wire I13868B;
wire I13258B;
wire I13259B;
wire g3261B;
wire I16074B;
wire I5136B;
wire I5137B;
wire I5460B;
wire I5461B;
wire I8605B;
wire I6770B;
wire I17401B;
wire g11449B;
wire g11448B;
wire g10231B;
wire I15716B;
wire I15717B;
wire I14210B;
wire I17567B;
wire I17569B;
wire I13876B;
wire I13878B;
wire I5606B;
wire I14442B;
wire I11996B;
wire I11997B;
wire I14277B;
wire I17568B;
wire I7321B;
wire I6990B;
wire g8847B;
wire I9006B;
wire I4985B;
wire I8651B;
wire I13544B;
wire I13545B;
wire I13894B;
wire I13895B;
wire I6136B;
wire I6138B;
wire I13076B;
wire g2205B;
wire I13260B;
wire I5501B;
wire I17586B;
wire I13900B;
wire I6201B;
wire g8826B;
wire I14216B;
wire I14217B;
wire I9007B;
wire I13559B;
wire I13561B;
wire g10229B;
wire I17492B;
wire I17493B;
wire I12214B;
wire I12215B;
wire I11262B;
wire I11263B;
wire I6225B;
wire I6226B;
wire I13307B;
wire I13309B;
wire I5676B;
wire I5677B;
wire I6826B;
wire I6827B;
wire g8190B;
wire I13308B;
wire I5879B;
wire I5880B;
wire g2792B;
wire g3061B;
wire I17585B;
wire I6881B;
wire I12138B;
wire g4605B;
wire I8728B;
wire I8729B;
wire I15871B;
wire I5866B;
wire I5867B;
wire I6793B;
wire I6487B;
wire I16080B;
wire I13893B;
wire I12115B;
wire I6748B;
wire I6224B;
wire I8805B;
wire I15878B;
wire I15880B;
wire I16030B;
wire I16031B;
wire I14271B;
wire I13267B;
wire I15616B;
wire I15617B;
wire I4964B;
wire I4966B;
wire I8752B;
wire I15432B;
wire g10438B;
wire g6032B;
wire g3011B;
wire I8480B;
wire I16086B;
wire I16087B;
wire g3734B;
wire I14218B;
wire I4955B;
wire g4639B;
wire I8786B;
wire g10480B;
wire I11914B;
wire I11915B;
wire g4619B;
wire I8770B;
wire I5516B;
wire g8541B;
wire I6188B;
wire I5891B;
wire I5892B;
wire I13766B;
wire I13767B;
wire I15258B;
wire I13266B;
wire I6825B;
wire I17283B;
wire g5277B;
wire I5035B;
wire g10359B;
wire I15879B;
wire I12114B;
wire I12107B;
wire g2500B;
wire g10430B;
wire g5999B;
wire I13285B;
wire I13877B;
wire I5893B;
wire g2795B;
wire I13560B;
wire g4259B;
wire I5166B;
wire I14614B;
wire I4965B;
wire I4943B;
wire I16023B;
wire I16059B;
wire g8737B;
wire I9576B;
wire I16052B;
wire I16053B;
wire I12004B;
wire g5573B;
wire I6837B;
wire I8730B;
wire I4978B;
wire I6177B;
wire I17051B;
wire I7864B;
wire I7865B;
wire I6665B;
wire I12216B;
wire I13554B;
wire I13284B;
wire I6137B;
wire I5529B;
wire I5530B;
wire I17282B;
wire I5618B;
wire I8662B;
wire I8664B;
wire I11916B;
wire g7717B;
wire I4971B;
wire I4972B;
wire I13273B;
wire I10509B;
wire I10508B;
wire I6778B;
wire I6779B;
wire I5469B;
wire g4251B;
wire I13546B;
wire I4996B;
wire I4997B;
wire I13539B;
wire I16032B;
wire I5323B;
wire I13538B;
wire I5540B;
wire I8778B;
wire g4286B;
wire I17052B;
wire I17053B;
wire I15898B;
wire g7978B;
wire g4227B;
wire I8561B;
wire I8762B;
wire I8751B;
wire I15907B;
wire I4973B;
wire I16024B;
wire I16025B;
wire g4455B;
wire I5341B;
wire I5342B;
wire I12137B;
wire I16088B;
wire g10483B;
wire I17289B;
wire g4630B;
wire I15609B;
wire I15608B;
wire g10436B;
wire g6023B;
wire I17459B;
wire I13301B;
wire I11981B;
wire I8663B;
wire I15718B;
wire I5284B;
wire g4607B;
wire g8840B;
wire g10441B;
wire g5345B;
wire g10432B;
wire g5938B;
wire I12021B;
wire I6489B;
wire I5528B;
wire I13659B;
wire I5343B;
wire I12039B;
wire I9008B;
wire I6488B;
wire I13888B;
wire I17494B;
wire I7684B;
wire g3221B;
wire I6324B;
wire I8590B;
wire I11243B;
wire g1737B;
wire g10324B;
wire g10239B;
wire g4974B;
wire g10322B;
wire g1736B;
wire g1955B;
wire g1956B;
wire g113B;
wire g1360B;
wire g1217B;
wire g755B;
wire g875B;
wire g1356B;
wire g874B;
wire FE_OFN370_g4525C;
wire FE_OFN369_g4525C;
wire FE_OFN368_g4525C;
wire FE_OFN367_g3521C;
wire FE_OFN366_g3521C;
wire FE_OFN365_g5361C;
wire FE_OFN364_g3015C;
wire FE_OFN363_I5565C;
wire FE_OFN362_g4525C;
wire FE_OFN360_g4525C;
wire FE_OFN359_g18C;
wire FE_OFN358_g3521C;
wire FE_OFN357_g3521C;
wire FE_OFN356_g5361C;
wire FE_OFN354_g5361C;
wire FE_OFN353_g5117C;
wire FE_OFN352_g109C;
wire FE_OFN351_g3913C;
wire FE_OFN350_g3121C;
wire FE_OFN349_I6424C;
wire FE_OFN348_g3015C;
wire FE_OFN347_g3914C;
wire FE_OFN346_g4381C;
wire FE_OFN345_g3015C;
wire FE_OFN344_g3586C;
wire FE_OFN343_I5565C;
wire FE_OFN340_I5565C;
wire FE_OFN339_g4525C;
wire FE_OFN337_g4525C;
wire FE_OFN336_g1690C;
wire FE_OFN335_g4737C;
wire FE_OFN334_g7045C;
wire FE_OFN333_g4294C;
wire FE_OFN332_g8748C;
wire FE_OFN331_g8696C;
wire FE_OFN330_g7638C;
wire FE_OFN329_g8763C;
wire FE_OFN328_g8709C;
wire FE_OFN325_g18C;
wire FE_OFN324_g18C;
wire FE_OFN322_g4449C;
wire FE_OFN321_g5261C;
wire FE_OFN320_g5361C;
wire FE_OFN319_g5361C;
wire FE_OFN318_g5361C;
wire FE_OFN316_g5361C;
wire FE_OFN315_g5117C;
wire FE_OFN312_g5117C;
wire FE_OFN310_g4336C;
wire FE_OFN308_I6424C;
wire FE_OFN307_g4010C;
wire FE_OFN306_g5128C;
wire FE_OFN305_g5151C;
wire FE_OFN304_g5151C;
wire FE_OFN303_g4678C;
wire FE_OFN302_g3913C;
wire FE_OFN300_g4002C;
wire FE_OFN299_g4457C;
wire FE_OFN298_g3015C;
wire FE_OFN297_g3015C;
wire FE_OFN296_g3914C;
wire FE_OFN294_g3914C;
wire FE_OFN293_g3015C;
wire FE_OFN292_g3015C;
wire FE_OFN291_g4880C;
wire FE_OFN290_g4880C;
wire FE_OFN289_g4679C;
wire FE_OFN288_g4263C;
wire FE_OFN287_g3586C;
wire FE_OFN284_g3586C;
wire FE_OFN283_I8869C;
wire FE_OFN282_g6165C;
wire FE_OFN281_g2216C;
wire FE_OFN280_g9536C;
wire FE_OFN279_g11157C;
wire FE_OFN278_g10927C;
wire FE_OFN277_g48C;
wire FE_OFN276_g48C;
wire FE_OFN275_g48C;
wire FE_OFN273_g85C;
wire FE_OFN271_g85C;
wire FE_OFN269_g109C;
wire FE_OFN267_g109C;
wire FE_OFN266_g18C;
wire FE_OFN260_g18C;
wire FE_OFN254_g461C;
wire FE_OFN253_g1786C;
wire FE_OFN252_g1791C;
wire FE_OFN251_g1801C;
wire FE_OFN250_g471C;
wire FE_OFN248_g466C;
wire FE_OFN247_g1771C;
wire FE_OFN245_g1690C;
wire FE_OFN241_g1690C;
wire FE_OFN240_g1110C;
wire FE_OFN239_g1796C;
wire FE_OFN238_g1781C;
wire FE_OFN237_g1806C;
wire FE_OFN236_g1776C;
wire FE_OFN235_g2024C;
wire FE_OFN234_g2024C;
wire FE_OFN233_I5565C;
wire FE_OFN230_I5565C;
wire FE_OFN229_g3880C;
wire FE_OFN227_g3880C;
wire FE_OFN226_g3880C;
wire FE_OFN225_g2276C;
wire FE_OFN224_g2276C;
wire FE_OFN223_g4401C;
wire FE_OFN221_g3440C;
wire FE_OFN219_g5557C;
wire FE_OFN218_g5557C;
wire FE_OFN217_g5013C;
wire FE_OFN213_g6003C;
wire FE_OFN211_g7246C;
wire FE_OFN210_g7246C;
wire FE_OFN209_g6863C;
wire FE_OFN207_g6863C;
wire FE_OFN206_g6863C;
wire FE_OFN204_g3664C;
wire FE_OFN200_g4921C;
wire FE_OFN199_g7697C;
wire FE_OFN198_g7697C;
wire FE_OFN196_g7697C;
wire FE_OFN195_g6488C;
wire FE_OFN192_g6488C;
wire FE_OFN191_g6488C;
wire FE_OFN189_g7638C;
wire FE_OFN187_g7638C;
wire FE_OFN184_I7048C;
wire FE_OFN180_g5354C;
wire FE_OFN179_g5354C;
wire FE_OFN178_g5354C;
wire FE_OFN177_g5919C;
wire FE_OFN176_g5151C;
wire FE_OFN168_g5361C;
wire FE_OFN166_g5361C;
wire FE_OFN164_g5361C;
wire FE_OFN161_g5361C;
wire FE_OFN160_I6424C;
wire FE_OFN155_g3121C;
wire FE_OFN154_g4640C;
wire FE_OFN153_g4640C;
wire FE_OFN147_g4682C;
wire FE_OFN146_g4682C;
wire FE_OFN144_g4682C;
wire FE_OFN142_g4682C;
wire FE_OFN141_g3829C;
wire FE_OFN137_g3829C;
wire FE_OFN136_g3863C;
wire FE_OFN134_g3863C;
wire FE_OFN133_g3015C;
wire FE_OFN132_g3015C;
wire FE_OFN131_g3015C;
wire FE_OFN119_g3015C;
wire FE_OFN118_g4807C;
wire FE_OFN117_g4807C;
wire FE_OFN116_g4807C;
wire FE_OFN115_g4807C;
wire FE_OFN113_g3914C;
wire FE_OFN111_g3914C;
wire FE_OFN110_g3586C;
wire FE_OFN103_g3586C;
wire FE_OFN102_g3586C;
wire FE_OFN100_g4421C;
wire FE_OFN99_g4421C;
wire FE_OFN97_I8869C;
wire FE_OFN96_g2169C;
wire FE_OFN95_g2216C;
wire FE_OFN93_g2216C;
wire FE_OFN92_g2216C;
wire FE_OFN91_g2172C;
wire FE_OFN90_I11360C;
wire FE_OFN89_I11360C;
wire FE_OFN88_g2178C;
wire FE_OFN87_g2176C;
wire FE_OFN86_g2176C;
wire FE_OFN85_g2176C;
wire FE_OFN84_g2176C;
wire FE_OFN83_g2176C;
wire FE_OFN82_g2176C;
wire FE_OFN81_g2176C;
wire FE_OFN80_g2175C;
wire FE_OFN79_g8700C;
wire FE_OFN76_g8700C;
wire FE_OFN73_g8858C;
wire FE_OFN72_g9292C;
wire FE_OFN71_g9292C;
wire FE_OFN70_g9490C;
wire FE_OFN69_g9392C;
wire FE_OFN68_g9392C;
wire FE_OFN67_g9367C;
wire FE_OFN64_g9536C;
wire FE_OFN63_g9474C;
wire FE_OFN62_g9274C;
wire FE_OFN61_g9624C;
wire FE_OFN60_g9624C;
wire FE_OFN59_g9432C;
wire FE_OFN57_g9432C;
wire FE_OFN56_g9052C;
wire FE_OFN54_g9052C;
wire FE_OFN53_g9173C;
wire FE_OFN52_g9173C;
wire FE_OFN51_g9111C;
wire FE_OFN50_g9030C;
wire FE_OFN49_g9030C;
wire FE_OFN48_g9151C;
wire FE_OFN47_g9151C;
wire FE_OFN46_g9125C;
wire FE_OFN45_g9125C;
wire FE_OFN44_g9125C;
wire FE_OFN42_g9205C;
wire FE_OFN40_g9240C;
wire FE_OFN39_g9223C;
wire FE_OFN35_g9785C;
wire FE_OFN34_g9785C;
wire FE_OFN33_g9454C;
wire FE_OFN32_g9454C;
wire FE_OFN27_g11519C;
wire FE_OFN21_g10702C;
wire FE_OFN20_g10702C;
wire FE_OFN18_g10702C;
wire FE_OFN17_g10702C;
wire FE_OFN15_g10702C;
wire FE_OFN14_g10702C;
wire FE_OFN13_g10702C;
wire FE_OFN10_g10702C;
wire FE_OFN9_g10702C;
wire FE_OFN8_g10702C;
wire FE_OFN7_g10702C;
wire FE_OFN4_g10950C;
wire FE_OFN3_g10950C;
wire FE_OFN0_g10950C;
wire g4500C;
wire g5529C;
wire g9968C;
wire g4682C;
wire g1707C;
wire g2299C;
wire g9291C;
wire g2807C;
wire I7048C;
wire g4130C;
wire g5024C;
wire g4338C;
wire g11596C;
wire g8147C;
wire g6551C;
wire g10865C;
wire g650C;
wire g1981C;
wire g8054C;
wire g3982C;
wire g9974C;
wire g1216C;
wire g546C;
wire g798C;
wire g3629C;
wire g7709C;
wire g8465C;
wire g8617C;
wire g4940C;
wire g4640C;
wire g135C;
wire g2078C;
wire g4565C;
wire g1918C;
wire g2340C;
wire g7684C;
wire g11519C;
wire g5935C;
wire g3800C;
wire g4736C;
wire g6941C;
wire g201C;
wire g2435C;
wire g4010C;
wire g1371C;
wire g2082C;
wire g4811C;
wire g5519C;
wire g49C;
wire g560C;
wire g6481C;
wire g6215C;
wire g10563C;
wire g10668C;
wire g70C;
wire g5013C;
wire g11221C;
wire g9508C;
wire g5212C;
wire g6529C;
wire g8709C;
wire g115C;
wire g2214C;
wire g5008C;
wire g3829C;
wire g9995C;
wire g10707C;
wire g3435C;
wire I7847C;
wire g5576C;
wire I13400C;
wire I5002C;
wire g10013C;
wire g10385C;
wire g9432C;
wire g3753C;
wire g4566C;
wire g254C;
wire I14326C;
wire g4722C;
wire g3348C;
wire g9696C;
wire g10408C;
wire I15968C;
wire g756C;
wire g818C;
wire g10937C;
wire g11060C;
wire g7242C;
wire g10336C;
wire I15855C;
wire g5229C;
wire g8940C;
wire g259C;
wire g10584C;
wire g10679C;
wire g4560C;
wire g10855C;
wire g369C;
wire g1968C;
wire I15503C;
wire g7996C;
wire g8110C;
wire g186C;
wire g2556C;
wire g3586C;
wire g10496C;
wire g3399C;
wire I7817C;
wire g158C;
wire g2222C;
wire g6907C;
wire g8226C;
wire I13373C;
wire g5405C;
wire I9880C;
wire g6155C;
wire g7246C;
wire g6638C;
wire g11647C;
wire g2744C;
wire g4094C;
wire g32C;
wire g3374C;
wire g4567C;
wire g8814C;
wire I14312C;
wire g10950C;
wire g9490C;
wire g11111C;
wire g4776C;
wire g5477C;
wire g6910C;
wire g10417C;
wire I15986C;
wire g713C;
wire g2237C;
wire g6488C;
wire g7712C;
wire g7897C;
wire g6828C;
wire g7638C;
wire g3015C;
wire g3121C;
wire I4917C;
wire g10800C;
wire g4300C;
wire g5420C;
wire g8019C;
wire I15956C;
wire g1840C;
wire g2557C;
wire g105C;
wire g9097C;
wire g6821C;
wire g3938C;
wire I5245C;
wire g253C;
wire g7682C;
wire g8267C;
wire g11478C;
wire g3698C;
wire g4379C;
wire g4144C;
wire g584C;
wire g131C;
wire g2254C;
wire g4289C;
wire g3992C;
wire g4777C;
wire I5424C;
wire g1776C;
wire g4585C;
wire g7934C;
wire g8089C;
wire g243C;
wire g2438C;
wire g6516C;
wire g8244C;
wire g4271C;
wire g4753C;
wire g8631C;
wire g4807C;
wire g10793C;
wire g7045C;
wire g5910C;
wire g9454C;
wire g686C;
wire g2212C;
wire I14299C;
wire g2563C;
wire g3141C;
wire g2478C;
wire g569C;
wire g35C;
wire g3215C;
wire g3710C;
wire I16252C;
wire g10726C;
wire g7516C;
wire g7920C;
wire g6824C;
wire g162C;
wire g2229C;
wire g9931C;
wire I15157C;
wire g11157C;
wire I15365C;
wire g79C;
wire I9279C;
wire g5361C;
wire g10558C;
wire g5248C;
wire g3880C;
wire g5557C;
wire g2172C;
wire g6759C;
wire g6502C;
wire g10797C;
wire g8241C;
wire I5044C;
wire g7685C;
wire g4471C;
wire g10780C;
wire g11625C;
wire g11372C;
wire g10007C;
wire I15287C;
wire g10771C;
wire I15290C;
wire g9720C;
wire g127C;
wire g2249C;
wire g5803C;
wire g11231C;
wire g11580C;
wire g5478C;
wire g11243C;
wire g4998C;
wire g10019C;
wire I5414C;
wire g4114C;
wire g11293C;
wire g2176C;
wire g4779C;
wire g5820C;
wire g8173C;
wire g3111C;
wire g3628C;
wire g4977C;
wire g6081C;
wire g255C;
wire g6533C;
wire I8503C;
wire g7460C;
wire g7910C;
wire g1984C;
wire g3688C;
wire g4285C;
wire g5867C;
wire g6354C;
wire g1690C;
wire g2031C;
wire g1857C;
wire I5510C;
wire g10405C;
wire g7932C;
wire g8085C;
wire g928C;
wire g7883C;
wire g10448C;
wire g5001C;
wire g8245C;
wire g3440C;
wire g4737C;
wire g8451C;
wire g8214C;
wire I13351C;
wire g3041C;
wire g10767C;
wire g10599C;
wire g10501C;
wire g3546C;
wire g8512C;
wire g2276C;
wire g6000C;
wire g6863C;
wire g10809C;
wire g10883C;
wire g5521C;
wire I14323C;
wire g11492C;
wire g932C;
wire g37C;
wire I6260C;
wire I9311C;
wire g4490C;
wire g8488C;
wire I5579C;
wire I9268C;
wire g4903C;
wire g10720C;
wire g10334C;
wire g10439C;
wire g6934C;
wire g5309C;
wire g5878C;
wire g4273C;
wire g7622C;
wire g6123C;
wire g7467C;
wire g774C;
wire g1990C;
wire g2248C;
wire g6838C;
wire g2045C;
wire g4905C;
wire g10798C;
wire g10785C;
wire g8187C;
wire I13436C;
wire g605C;
wire g2399C;
wire g7204C;
wire g6830C;
wire g6716C;
wire g8944C;
wire I5254C;
wire g5543C;
wire I5410C;
wire g5300C;
wire g8921C;
wire g8745C;
wire g8849C;
wire g6096C;
wire I7752C;
wire g6003C;
wire g3431C;
wire I7840C;
wire g10852C;
wire g6733C;
wire g7562C;
wire g6548C;
wire g1419C;
wire I9810C;
wire g5502C;
wire g260C;
wire g4679C;
wire g6823C;
wire g4890C;
wire g7981C;
wire g2579C;
wire g3776C;
wire g572C;
wire g3381C;
wire g10863C;
wire g971C;
wire g2008C;
wire g8039C;
wire g6526C;
wire g1900C;
wire g2336C;
wire g10664C;
wire g7189C;
wire g5278C;
wire g8923C;
wire g5173C;
wire g3521C;
wire I14306C;
wire g10712C;
wire I9296C;
wire g4264C;
wire g2178C;
wire g6755C;
wire g2791C;
wire I6962C;
wire g5226C;
wire g704C;
wire g2230C;
wire g4437C;
wire g11514C;
wire g7505C;
wire g38C;
wire g9507C;
wire g10411C;
wire I15974C;
wire g4506C;
wire g1834C;
wire g2550C;
wire g10348C;
wire g10400C;
wire I9282C;
wire I5584C;
wire g9324C;
wire g3664C;
wire g10001C;
wire g5526C;
wire g7697C;
wire g231C;
wire g2395C;
wire I5395C;
wire g4788C;
wire g4465C;
wire g8289C;
wire g6403C;
wire g8203C;
wire I15510C;
wire g5403C;
wire g6902C;
wire g6015C;
wire g11340C;
wire g6542C;
wire I5406C;
wire g3744C;
wire g581C;
wire I4883C;
wire g4537C;
wire g7688C;
wire g882C;
wire g2481C;
wire g6507C;
wire g10485C;
wire I4935C;
wire g10683C;
wire I9308C;
wire I5070C;
wire g5556C;
wire g8505C;
wire g8603C;
wire g11641C;
wire g3423C;
wire g4787C;
wire I9332C;
wire g10765C;
wire g6447C;
wire g4801C;
wire g11305C;
wire g3092C;
wire g6126C;
wire g4281C;
wire g5493C;
wire g5613C;
wire g639C;
wire g10414C;
wire g7986C;
wire g8255C;
wire g8000C;
wire g8081C;
wire g814C;
wire I9479C;
wire I4780C;
wire g2216C;
wire g10522C;
wire I5383C;
wire g8060C;
wire g7191C;
wire g8746C;
wire g8783C;
wire g10557C;
wire g5150C;
wire I5445C;
wire g4449C;
wire I4866C;
wire g6469C;
wire g7696C;
wire g10452C;
wire g4498C;
wire g8744C;
wire g8828C;
wire g2034C;
wire g2677C;
wire g5514C;
wire g6627C;
wire g4893C;
wire g10268C;
wire g10361C;
wire g3737C;
wire g9257C;
wire g9525C;
wire g5194C;
wire g668C;
wire g2198C;
wire g3418C;
wire I7771C;
wire g6901C;
wire g8043C;
wire g5263C;
wire g6929C;
wire g5857C;
wire g3523C;
wire g8049C;
wire g4529C;
wire g9699C;
wire g722C;
wire g2241C;
wire g6786C;
wire g7218C;
wire g7681C;
wire g6234C;
wire g5824C;
wire g7101C;
wire g10864C;
wire g7651C;
wire g7914C;
wire g986C;
wire I13427C;
wire g8816C;
wire I14319C;
wire I5430C;
wire g2175C;
wire g10862C;
wire I15980C;
wire g11077C;
wire I9259C;
wire g7683C;
wire I16717C;
wire I5388C;
wire I9326C;
wire g153C;
wire g2211C;
wire g3222C;
wire g3983C;
wire g4678C;
wire g3101C;
wire g3543C;
wire I5053C;
wire g9268C;
wire g5942C;
wire g10331C;
wire g10421C;
wire g10721C;
wire g8051C;
wire g2118C;
wire g10383C;
wire g6541C;
wire g936C;
wire g9088C;
wire g139C;
wire g2083C;
wire I6360C;
wire g10773C;
wire g8193C;
wire I4992C;
wire g6523C;
wire I16982C;
wire g8546C;
wire g8599C;
wire g794C;
wire g1828C;
wire g2061C;
wire g746C;
wire g2187C;
wire I9383C;
wire g5404C;
wire g11393C;
wire g5258C;
wire g1845C;
wire g2271C;
wire g1400C;
wire g2446C;
wire g8265C;
wire g2984C;
wire g11561C;
wire g11575C;
wire g822C;
wire g4765C;
wire g4334C;
wire g1936C;
wire g2345C;
wire g11233C;
wire g7950C;
wire g8106C;
wire g6586C;
wire g6908C;
wire g8768C;
wire g8885C;
wire g563C;
wire g33C;
wire g5808C;
wire I5418C;
wire g1361C;
wire g2016C;
wire g5271C;
wire g6333C;
wire g10515C;
wire g7692C;
wire I9273C;
wire g6045C;
wire g123C;
wire g731C;
wire g2251C;
wire g1988C;
wire g2047C;
wire g10927C;
wire g7590C;
wire g2275C;
wire g6468C;
wire g10782C;
wire g10886C;
wire g6672C;
wire g6840C;
wire g5230C;
wire g549C;
wire g8743C;
wire g8858C;
wire g3354C;
wire g4671C;
wire g5914C;
wire g7705C;
wire g7953C;
wire g8115C;
wire g10025C;
wire g1218C;
wire g2017C;
wire I5101C;
wire g6038C;
wire g1882C;
wire g2328C;
wire I5057C;
wire g1868C;
wire g2542C;
wire g4488C;
wire g1891C;
wire g2330C;
wire g3863C;
wire g6471C;
wire g11303C;
wire I9276C;
wire g7949C;
wire I5041C;
wire g782C;
wire g1992C;
wire I5441C;
wire g1110C;
wire g4365C;
wire g5266C;
wire g8234C;
wire I13364C;
wire g4158C;
wire g10663C;
wire g8920C;
wire g4283C;
wire I4859C;
wire g10788C;
wire g1397C;
wire g2456C;
wire g7512C;
wire g7919C;
wire g4484C;
wire I17413C;
wire I9346C;
wire g643C;
wire g1976C;
wire g7952C;
wire g865C;
wire I4820C;
wire I5435C;
wire g8815C;
wire I14315C;
wire g3008C;
wire g4467C;
wire g9713C;
wire g4290C;
wire g7527C;
wire g4770C;
wire g9474C;
wire g36C;
wire g5842C;
wire I9265C;
wire g7671C;
wire g8056C;
wire g8700C;
wire g4381C;
wire g5396C;
wire g1854C;
wire g7203C;
wire I6273C;
wire g10382C;
wire g10583C;
wire g10629C;
wire g8045C;
wire g7843C;
wire g2652C;
wire g754C;
wire g2057C;
wire g3539C;
wire g4263C;
wire g8269C;
wire I9349C;
wire I13323C;
wire g1386C;
wire g2549C;
wire g5261C;
wire g3104C;
wire g3419C;
wire g3425C;
wire I7829C;
wire g9802C;
wire g806C;
wire g6537C;
wire I13338C;
wire g5221C;
wire g3086C;
wire g2253C;
wire g4902C;
wire g6080C;
wire I9371C;
wire g5485C;
wire g6059C;
wire g4089C;
wire I5588C;
wire g7664C;
wire g7907C;
wire g4673C;
wire g8551C;
wire g5126C;
wire g10866C;
wire g10597C;
wire g11603C;
wire g6332C;
wire g4231C;
wire g9526C;
wire g207C;
wire g2570C;
wire g7473C;
wire g7915C;
wire I4783C;
wire g1991C;
wire g7677C;
wire g64C;
wire g11249C;
wire g636C;
wire g2506C;
wire g11348C;
wire g10779C;
wire g11488C;
wire g3491C;
wire g40C;
wire g3438C;
wire I7852C;
wire g757C;
wire g5354C;
wire g5295C;
wire g5918C;
wire g6894C;
wire g3513C;
wire g1713C;
wire I6240C;
wire g258C;
wire g591C;
wire g2374C;
wire g9424C;
wire g4076C;
wire g6534C;
wire g58C;
wire g3793C;
wire g6928C;
wire g7686C;
wire g3414C;
wire I7825C;
wire g8055C;
wire g11291C;
wire g237C;
wire g2420C;
wire g3209C;
wire g4739C;
wire g5509C;
wire g6833C;
wire g1958C;
wire g6918C;
wire g4608C;
wire I4948C;
wire g6915C;
wire g6911C;
wire I5060C;
wire g8812C;
wire I9237C;
wire g4553C;
wire g7441C;
wire g5996C;
wire g8047C;
wire g1786C;
wire g6653C;
wire g7438C;
wire g6832C;
wire I5047C;
wire g4771C;
wire g11481C;
wire g10857C;
wire g7947C;
wire g8100C;
wire g3681C;
wire g7918C;
wire I5427C;
wire g6478C;
wire g4117C;
wire g6897C;
wire g6042C;
wire I9717C;
wire g119C;
wire g11229C;
wire g1453C;
wire g2410C;
wire g10402C;
wire g4342C;
wire g4330C;
wire g8221C;
wire g1927C;
wire g2343C;
wire g11609C;
wire g10859C;
wire g6054C;
wire g6508C;
wire g6531C;
wire g8050C;
wire g8261C;
wire I9290C;
wire g11376C;
wire g580C;
wire I4876C;
wire g802C;
wire g8559C;
wire I9769C;
wire g2260C;
wire g10556C;
wire g148C;
wire g2202C;
wire g7032C;
wire g8390C;
wire g8548C;
wire g590C;
wire g2518C;
wire g4548C;
wire g4293C;
wire I16507C;
wire g5390C;
wire g4561C;
wire g8233C;
wire g1289C;
wire g8200C;
wire g4294C;
wire g76C;
wire g8767C;
wire g3071C;
wire g3723C;
wire I15962C;
wire g940C;
wire g7987C;
wire g8094C;
wire g1861C;
wire g2050C;
wire g1987C;
wire g4480C;
wire g11483C;
wire g1351C;
wire g10702C;
wire g5863C;
wire g2273C;
wire g5392C;
wire g9082C;
wire g5838C;
wire g8270C;
wire g10776C;
wire g2024C;
wire g2777C;
wire g6513C;
wire g9272C;
wire g10732C;
wire g1411C;
wire g10898C;
wire g869C;
wire g8052C;
wire g4325C;
wire g3368C;
wire g762C;
wire g4421C;
wire I8869C;
wire g5319C;
wire g8766C;
wire g10555C;
wire g586C;
wire g61C;
wire g6205C;
wire g778C;
wire g622C;
wire g8820C;
wire I9329C;
wire g11199C;
wire g9124C;
wire g6839C;
wire g6522C;
wire g10936C;
wire g7852C;
wire g7923C;
wire g11320C;
wire g6841C;
wire g10328C;
wire g10431C;
wire g8769C;
wire g6224C;
wire g2208C;
wire g11349C;
wire g4782C;
wire g6470C;
wire g11225C;
wire g5755C;
wire g4292C;
wire g1212C;
wire g6515C;
wire g3003C;
wire g3760C;
wire g9710C;
wire g5117C;
wire g3631C;
wire g5182C;
wire g11430C;
wire I9368C;
wire g10791C;
wire g5004C;
wire g1806C;
wire g7632C;
wire g11485C;
wire I5399C;
wire g6331C;
wire g1718C;
wire g2424C;
wire g5257C;
wire g8053C;
wire g4518C;
wire g7550C;
wire g219C;
wire g2077C;
wire g3103C;
wire g4764C;
wire g7913C;
wire g1989C;
wire g3068C;
wire g6109C;
wire I15500C;
wire g5763C;
wire g6480C;
wire g6795C;
wire g6449C;
wire g8194C;
wire g2257C;
wire g5201C;
wire g5269C;
wire g7497C;
wire g876C;
wire g2444C;
wire g1107C;
wire g8938C;
wire g7990C;
wire g8099C;
wire g4238C;
wire g8775C;
wire g4891C;
wire g8266C;
wire g11290C;
wire g6501C;
wire g10570C;
wire g10676C;
wire g6334C;
wire g786C;
wire g1993C;
wire g10719C;
wire g1104C;
wire g4727C;
wire g4274C;
wire g8765C;
wire g6916C;
wire g8811C;
wire I14303C;
wire g5174C;
wire I5525C;
wire I14330C;
wire g583C;
wire I4900C;
wire g11308C;
wire g3060C;
wire g5847C;
wire g10554C;
wire g10784C;
wire g2979C;
wire g599C;
wire g2382C;
wire g7680C;
wire g10396C;
wire g3784C;
wire g11425C;
wire I14295C;
wire g1346C;
wire I9293C;
wire I5815C;
wire g4002C;
wire g7062C;
wire g3479C;
wire g5548C;
wire g6131C;
wire g2449C;
wire g6820C;
wire g3390C;
wire g5627C;
wire g3501C;
wire g4340C;
wire I13385C;
wire g143C;
wire g2095C;
wire g1771C;
wire g257C;
wire g2297C;
wire g262C;
wire g6922C;
wire g1969C;
wire g6747C;
wire g11391C;
wire g8818C;
wire g8649C;
wire g9555C;
wire g6071C;
wire g1796C;
wire g7942C;
wire g8095C;
wire g6718C;
wire g611C;
wire g2364C;
wire g10858C;
wire g55C;
wire g1864C;
wire g2054C;
wire g2018C;
wire g2725C;
wire g627C;
wire g8926C;
wire g4239C;
wire g11602C;
wire g8041C;
wire g5503C;
wire g646C;
wire g1980C;
wire g981C;
wire g8164C;
wire g883C;
wire I6220C;
wire g582C;
wire I4891C;
wire g8922C;
wire g5536C;
wire g578C;
wire g5810C;
wire g7067C;
wire g8236C;
wire g11605C;
wire g8048C;
wire g6528C;
wire g1909C;
wire g2338C;
wire g34C;
wire g6524C;
wire g7446C;
wire g3056C;
wire g3475C;
wire g7258C;
wire g7219C;
wire g8046C;
wire g3706C;
wire g4822C;
wire g11482C;
wire g10381C;
wire g4477C;
wire g10333C;
wire g10437C;
wire g4456C;
wire g2310C;
wire g3039C;
wire g6923C;
wire g4255C;
wire g878C;
wire g790C;
wire g4732C;
wire g8937C;
wire g4752C;
wire g6538C;
wire g10339C;
wire g3524C;
wire g11306C;
wire g7183C;
wire g4778C;
wire g6165C;
wire g6895C;
wire g588C;
wire g11223C;
wire g6163C;
wire g6179C;
wire g9052C;
wire g9505C;
wire g9721C;
wire g654C;
wire g2268C;
wire g8776C;
wire g6827C;
wire g461C;
wire g4309C;
wire g9331C;
wire g7244C;
wire g7586C;
wire g7930C;
wire g5222C;
wire g11300C;
wire g10718C;
wire g213C;
wire g2070C;
wire g3906C;
wire g579C;
wire g5445C;
wire g11227C;
wire g6088C;
wire g658C;
wire g2331C;
wire g1365C;
wire g2406C;
wire g8206C;
wire I13332C;
wire g6679C;
wire g11636C;
wire g11239C;
wire g11219C;
wire g225C;
wire g2087C;
wire g2117C;
wire g2801C;
wire g3062C;
wire g3738C;
wire g9266C;
wire g9760C;
wire g11608C;
wire g8059C;
wire g8771C;
wire g2459C;
wire g6035C;
wire g1811C;
wire g7106C;
wire g471C;
wire g6198C;
wire g7992C;
wire g8105C;
wire g2169C;
wire g8973C;
wire g617C;
wire g2369C;
wire g6834C;
wire g197C;
wire g2407C;
wire g1962C;
wire g5148C;
wire I14642C;
wire g5836C;
wire g7134C;
wire I15514C;
wire g10795C;
wire g11083C;
wire g11276C;
wire g10770C;
wire g1810C;
wire g9271C;
wire g677C;
wire g2203C;
wire g587C;
wire I5497C;
wire I13421C;
wire g10494C;
wire g8773C;
wire g3462C;
wire I16220C;
wire g3662C;
wire g6740C;
wire g10484C;
wire g7143C;
wire g8939C;
wire g1703C;
wire g2028C;
wire g8772C;
wire g4336C;
wire g2067C;
wire g1814C;
wire g2564C;
wire g6093C;
wire g6500C;
wire g1407C;
wire g3705C;
wire g10500C;
wire g2794C;
wire g4065C;
wire g4243C;
wire g4934C;
wire g6485C;
wire g8777C;
wire g6244C;
wire g5304C;
wire g11640C;
wire g3814C;
wire g4784C;
wire g11487C;
wire g9110C;
wire g1822C;
wire g2571C;
wire g11380C;
wire g1950C;
wire g826C;
wire g9269C;
wire g7054C;
wire g1975C;
wire g7236C;
wire g2774C;
wire g3247C;
wire g3967C;
wire g11314C;
wire g585C;
wire g5276C;
wire g9150C;
wire g1389C;
wire g2396C;
wire g11298C;
wire g7202C;
wire g6819C;
wire g2987C;
wire g758C;
wire g11539C;
wire g1336C;
wire g108C;
wire g5317C;
wire g67C;
wire g10453C;
wire g6243C;
wire g6514C;
wire g8817C;
wire g8810C;
wire g1206C;
wire I6277C;
wire g1368C;
wire g2381C;
wire g9313C;
wire g10387C;
wire g6983C;
wire g8366C;
wire g8509C;
wire g7450C;
wire g7905C;
wire g4473C;
wire g6577C;
wire g1341C;
wire g1374C;
wire g2421C;
wire g3200C;
wire g4001C;
wire g8040C;
wire g5255C;
wire g6900C;
wire g8042C;
wire g11490C;
wire g11515C;
wire g8230C;
wire g6546C;
wire g3485C;
wire g1383C;
wire g2562C;
wire g6697C;
wire g8574C;
wire g5770C;
wire I11360C;
wire g8889C;
wire g10711C;
wire g9719C;
wire g11312C;
wire g5287C;
wire g11107C;
wire g1791C;
wire g6351C;
wire g9778C;
wire g6479C;
wire g3120C;
wire g3765C;
wire g5814C;
wire g5849C;
wire g1101C;
wire g575C;
wire g10559C;
wire g5219C;
wire g7240C;
wire I9352C;
wire g8819C;
wire g9256C;
wire g261C;
wire g6656C;
wire g976C;
wire g736C;
wire g1424C;
wire g1377C;
wire g2074C;
wire g6906C;
wire g10717C;
wire g4759C;
wire g5189C;
wire g8770C;
wire g6392C;
wire g6621C;
wire g11610C;
wire g4582C;
wire g6432C;
wire g7454C;
wire g7908C;
wire g8264C;
wire g11604C;
wire g9764C;
wire g2161C;
wire g3291C;
wire g7245C;
wire g2510C;
wire g256C;
wire g2439C;
wire g3207C;
wire g810C;
wire g11486C;
wire g12C;
wire g2126C;
wire g7581C;
wire g10799C;
wire I15507C;
wire I9221C;
wire g114C;
wire g1964C;
wire g10357C;
wire g6439C;
wire g8507C;
wire g8688C;
wire g7133C;
wire g8642C;
wire g8044C;
wire g8254C;
wire g11549C;
wire g1357C;
wire g2023C;
wire g7379C;
wire g11232C;
wire g11607C;
wire g6573C;
wire g3506C;
wire g3407C;
wire g770C;
wire g6193C;
wire g3108C;
wire g3408C;
wire g248C;
wire g2451C;
wire g7225C;
wire g8220C;
wire g7231C;
wire g4576C;
wire g3943C;
wire g4904C;
wire g8806C;
wire g11292C;
wire g6822C;
wire g7624C;
wire g3661C;
wire I15861C;
wire g73C;
wire g1801C;
wire g8327C;
wire g6912C;
wire g6898C;
wire g554C;
wire g8146C;
wire I5020C;
wire g5421C;
wire g1766C;
wire g7994C;
wire g8103C;
wire g1362C;
wire g2434C;
wire g3913C;
wire g6702C;
wire g4880C;
wire g8696C;
wire g868C;
wire g8813C;
wire I14309C;
wire g1945C;
wire g2347C;
wire g6924C;
wire g5308C;
wire g7574C;
wire g11310C;
wire g11294C;
wire g5852C;
wire g2970C;
wire g6026C;
wire g10369C;
wire g5286C;
wire g4554C;
wire g8024C;
wire g8945C;
wire g4804C;
wire g6525C;
wire g1380C;
wire g2060C;
wire g6019C;
wire g6617C;
wire g8210C;
wire g5083C;
wire g3585C;
wire g589C;
wire g7541C;
wire g4760C;
wire g26C;
wire g2479C;
wire g10860C;
wire g10502C;
wire g11579C;
wire g11639C;
wire g9814C;
wire g5030C;
wire g39C;
wire g6826C;
wire g2303C;
wire g9773C;
wire g52C;
wire g7626C;
wire g5200C;
wire g4457C;
wire g6829C;
wire g7211C;
wire g466C;
wire g456C;
wire g7660C;
wire g10722C;
wire g8887C;
wire g11484C;
wire g11286C;
wire g6002C;
wire g11606C;
wire g11217C;
wire g10454C;
wire g6757C;
wire g6216C;
wire g8941C;
wire g10856C;
wire g4892C;
wire g7903C;
wire g6930C;
wire g8250C;
wire g5250C;
wire g4525C;
wire g6049C;
wire g8943C;
wire g10861C;
wire g192C;
wire g2475C;
wire g8779C;
wire g766C;
wire g5484C;
wire g557C;
wire g11203C;
wire g3304C;
wire g6557C;
wire g4482C;
wire g1781C;
wire g5190C;
wire g6180C;
wire g5274C;
wire g8774C;
wire g10325C;
wire g10444C;
wire g566C;
wire g8260C;
wire g6099C;
wire g10401C;
wire g6831C;
wire g6068C;
wire g7137C;
wire g7917C;
wire g9473C;
wire g1965C;
wire g6545C;
wire g11547C;
wire g7257C;
wire g6909C;
wire g8384C;
wire g1872C;
wire g2503C;
wire g11392C;
wire g6506C;
wire g8883C;
wire g695C;
wire g2224C;
wire g6728C;
wire g10724C;
wire g4556C;
wire g3070C;
wire g2250C;
wire g11103C;
wire g9900C;
wire g845C;
wire g11095C;
wire g1645C;
wire g4973C;
wire g7389C;
wire g7465C;
wire g7888C;
wire g1642C;
wire g4969C;
wire g8224C;
wire g2892C;
wire g5686C;
wire g10308C;
wire g4123C;
wire g8120C;
wire g287C;
wire g6788C;
wire g4824C;
wire g5598C;
wire g278C;
wire g9694C;
wire g10495C;
wire g1684C;
wire g2945C;
wire g11190C;
wire g8639C;
wire g8789C;
wire g9728C;
wire g9563C;
wire g9852C;
wire g1053C;
wire g5625C;
wire g995C;
wire g4875C;
wire g1574C;
wire g9701C;
wire g7138C;
wire g10752C;
wire g11058C;
wire g11211C;
wire g435C;
wire g11024C;
wire g8307C;
wire g8547C;
wire g10669C;
wire g691C;
wire g7707C;
wire g3813C;
wire g4884C;
wire g4839C;
wire g1561C;
wire g9870C;
wire g6640C;
wire g9240C;
wire g9650C;
wire g5687C;
wire g7957C;
wire g3512C;
wire g7449C;
wire g1011C;
wire g4235C;
wire g345C;
wire g4343C;
wire g11296C;
wire g1C;
wire g9292C;
wire g9594C;
wire g1160C;
wire g9923C;
wire g9367C;
wire g9943C;
wire g1721C;
wire g5525C;
wire g440C;
wire g8876C;
wire g476C;
wire g10564C;
wire g10705C;
wire g9913C;
wire g9624C;
wire g9934C;
wire g6225C;
wire g1240C;
wire g6324C;
wire g10686C;
wire g1223C;
wire g6540C;
wire g8663C;
wire g1308C;
wire g11581C;
wire g6206C;
wire g452C;
wire g3989C;
wire g7260C;
wire g7730C;
wire g1235C;
wire g7504C;
wire g1887C;
wire g7185C;
wire I5689C;
wire I5690C;
wire g7881C;
wire g11070C;
wire g9736C;
wire g9859C;
wire g8877C;
wire g2274C;
wire g11590C;
wire g6199C;
wire g8932C;
wire g1730C;
wire g5545C;
wire g5180C;
wire g1615C;
wire g5591C;
wire g8412C;
wire g8556C;
wire g374C;
wire g11094C;
wire g5044C;
wire g5853C;
wire g6245C;
wire g4360C;
wire g8930C;
wire g5507C;
wire g3087C;
wire g11150C;
wire g8302C;
wire g8464C;
wire g272C;
wire g9692C;
wire g1428C;
wire g4996C;
wire g7131C;
wire g421C;
wire g11019C;
wire g9951C;
wire g9536C;
wire g9960C;
wire g11196C;
wire g11018C;
wire g10550C;
wire g10595C;
wire g10433C;
wire g10544C;
wire g10623C;
wire g4878C;
wire g4838C;
wire g5204C;
wire g8609C;
wire g8844C;
wire g6185C;
wire g6701C;
wire g10725C;
wire g5100C;
wire g1089C;
wire g4882C;
wire g8731C;
wire g1504C;
wire g5128C;
wire g1932C;
wire g6886C;
wire g8415C;
wire g8557C;
wire g8966C;
wire g8071C;
wire g11597C;
wire g9722C;
wire g9785C;
wire g9828C;
wire g1672C;
wire g2918C;
wire g9725C;
wire g9830C;
wire g8955C;
wire g4C;
wire g9592C;
wire g1618C;
wire g5123C;
wire g6078C;
wire g7059C;
wire g7459C;
wire g861C;
wire g11102C;
wire g709C;
wire g7718C;
wire g7535C;
wire g1577C;
wire g9703C;
wire g5528C;
wire g9911C;
wire g9932C;
wire g1636C;
wire g5530C;
wire g2760C;
wire g8629C;
wire g6187C;
wire g6887C;
wire g5605C;
wire g6228C;
wire g1275C;
wire g6322C;
wire I6337C;
wire I6338C;
wire g8967C;
wire g1458C;
wire g5010C;
wire g3275C;
wire g1678C;
wire g2895C;
wire g7721C;
wire g1549C;
wire g9866C;
wire g1534C;
wire g9716C;
wire g10744C;
wire g10808C;
wire g1231C;
wire g3047C;
wire g3685C;
wire g4492C;
wire g8614C;
wire g8822C;
wire g10560C;
wire g11456C;
wire g9724C;
wire g9848C;
wire g4714C;
wire g6550C;
wire g5172C;
wire g10642C;
wire g2531C;
wire g3284C;
wire g284C;
wire g302C;
wire g9855C;
wire g1630C;
wire g5618C;
wire g6891C;
wire g7940C;
wire g312C;
wire g11085C;
wire g396C;
wire g1432C;
wire g4968C;
wire g8646C;
wire g8837C;
wire g9125C;
wire g9644C;
wire g1546C;
wire g5804C;
wire g8300C;
wire g8462C;
wire I6330C;
wire g333C;
wire g11156C;
wire g293C;
wire g6342C;
wire g1552C;
wire g9867C;
wire g1537C;
wire g9717C;
wire g4871C;
wire g10435C;
wire g426C;
wire g7741C;
wire g1327C;
wire g9151C;
wire g9386C;
wire g8607C;
wire g8842C;
wire g8C;
wire g9599C;
wire g8974C;
wire g9274C;
wire g5518C;
wire g9111C;
wire g9614C;
wire g4122C;
wire g4610C;
wire g7217C;
wire g11557C;
wire g1675C;
wire g2911C;
wire g11210C;
wire g7466C;
wire g9918C;
wire g9939C;
wire g11279C;
wire g10513C;
wire g10440C;
wire I16145C;
wire g10518C;
wire g1129C;
wire g7055C;
wire g1095C;
wire g5264C;
wire g1265C;
wire g6329C;
wire g8176C;
wire g7510C;
wire g8005C;
wire g3281C;
wire g4099C;
wire g11601C;
wire g11187C;
wire g6746C;
wire g6221C;
wire g8630C;
wire g9622C;
wire g10923C;
wire g11143C;
wire g9886C;
wire g9676C;
wire g9904C;
wire g8733C;
wire g348C;
wire g6624C;
wire g530C;
wire g11169C;
wire g8073C;
wire g9706C;
wire g9512C;
wire g9841C;
wire g5592C;
wire g5882C;
wire g8645C;
wire g8796C;
wire g534C;
wire g11168C;
wire g1015C;
wire g4269C;
wire g727C;
wire g1047C;
wire g5611C;
wire g673C;
wire g8069C;
wire g1567C;
wire g9695C;
wire g10304C;
wire g8305C;
wire g8469C;
wire g1071C;
wire g4712C;
wire g5762C;
wire g6576C;
wire g10622C;
wire g5217C;
wire g11015C;
wire g5674C;
wire g9173C;
wire g9359C;
wire g8960C;
wire g9223C;
wire g11556C;
wire g1595C;
wire g9858C;
wire g5541C;
wire g363C;
wire g4534C;
wire g1499C;
wire g5897C;
wire g6177C;
wire g6699C;
wire g6855C;
wire g3098C;
wire g3804C;
wire g5680C;
wire g9642C;
wire g1528C;
wire g5744C;
wire g8399C;
wire g1762C;
wire g9030C;
wire g9447C;
wire g1849C;
wire g516C;
wire g11178C;
wire g8414C;
wire g8510C;
wire g1296C;
wire g6319C;
wire g11186C;
wire g1681C;
wire g2951C;
wire g6352C;
wire g9205C;
wire g9595C;
wire g4109C;
wire g4831C;
wire g1654C;
wire g5492C;
wire g8934C;
wire g10312C;
wire g6186C;
wire g9612C;
wire g1738C;
wire g9417C;
wire g9914C;
wire g9935C;
wire g10658C;
wire g10745C;
wire g956C;
wire g11216C;
wire g8971C;
wire g9328C;
wire g11587C;
wire g1245C;
wire g6325C;
wire g431C;
wire g7368C;
wire g552C;
wire g6083C;
wire g1227C;
wire g6544C;
wire g5476C;
wire g7743C;
wire g1083C;
wire g4869C;
wire g1598C;
wire g5722C;
wire g5813C;
wire g6790C;
wire g8408C;
wire g10761C;
wire g7734C;
wire g7926C;
wire g8136C;
wire g5569C;
wire g401C;
wire g9392C;
wire g9902C;
wire g8623C;
wire g1657C;
wire g5500C;
wire g2496C;
wire g3010C;
wire g5877C;
wire g6756C;
wire g8972C;
wire g336C;
wire g6622C;
wire g11612C;
wire g1311C;
wire g9366C;
wire g11230C;
wire g1284C;
wire g1215C;
wire g4364C;
wire g9649C;
wire g1543C;
wire g5795C;
wire g1524C;
wire g5737C;
wire g1753C;
wire g4054C;
wire g5823C;
wire g6345C;
wire g11275C;
wire g296C;
wire g9851C;
wire g5802C;
wire g6763C;
wire g416C;
wire g10511C;
wire g10509C;
wire g10507C;
wire I16142C;
wire g1571C;
wire g9698C;
wire g1032C;
wire g4725C;
wire g9954C;
wire g9964C;
wire g1663C;
wire g5523C;
wire g8402C;
wire g8550C;
wire g8611C;
wire g8845C;
wire g2081C;
wire g281C;
wire g6359C;
wire g1324C;
wire g11586C;
wire g5147C;
wire g11007C;
wire g5104C;
wire g4821C;
wire g5099C;
wire g5919C;
wire g1627C;
wire g5499C;
wire g3529C;
wire g4389C;
wire g3497C;
wire g6416C;
wire g1444C;
wire g4990C;
wire g9010C;
wire g9619C;
wire I6630C;
wire g6047C;
wire g953C;
wire g9652C;
wire g10505C;
wire g10469C;
wire g9711C;
wire g9519C;
wire g9843C;
wire g1074C;
wire g5273C;
wire g11465C;
wire g4348C;
wire g11237C;
wire g9731C;
wire g9834C;
wire g6654C;
wire g1041C;
wire g5444C;
wire g3714C;
wire g11285C;
wire g9598C;
wire g8097C;
wire g8726C;
wire g4816C;
wire g6880C;
wire g1157C;
wire g3287C;
wire g10759C;
wire g9917C;
wire g9938C;
wire g10652C;
wire g10758C;
wire g406C;
wire g9891C;
wire g9909C;
wire g6663C;
wire g7127C;
wire g11165C;
wire g1260C;
wire g6328C;
wire g8401C;
wire g5125C;
wire g11006C;
wire g1080C;
wire g4865C;
wire g1077C;
wire g4715C;
wire g2325C;
wire g4604C;
wire g5513C;
wire g965C;
wire g11222C;
wire g1145C;
wire g6554C;
wire g7732C;
wire g9586C;
wire g4401C;
wire g4104C;
wire g5178C;
wire g4584C;
wire g7472C;
wire g11253C;
wire g9860C;
wire g11600C;
wire g1586C;
wire g9645C;
wire g11236C;
wire g3106C;
wire g4162C;
wire g553C;
wire g6090C;
wire g269C;
wire g9691C;
wire g11316C;
wire g501C;
wire g11175C;
wire g664C;
wire g8068C;
wire g9607C;
wire g9952C;
wire g9962C;
wire g6348C;
wire g9659C;
wire g1318C;
wire g9358C;
wire I6316C;
wire I6317C;
wire g1711C;
wire g4486C;
wire g8995C;
wire g9587C;
wire g5632C;
wire g8965C;
wire g991C;
wire g4881C;
wire g11209C;
wire g8715C;
wire g8848C;
wire g3263C;
wire g4070C;
wire g6463C;
wire g1896C;
wire g7820C;
wire g448C;
wire g11021C;
wire g1044C;
wire g5917C;
wire g6619C;
wire g1300C;
wire g6318C;
wire g6872C;
wire g11201C;
wire g10489C;
wire g10514C;
wire g4006C;
wire g299C;
wire g9853C;
wire g11274C;
wire g8119C;
wire g1747C;
wire g9420C;
wire g5233C;
wire g7092C;
wire g6549C;
wire g11464C;
wire g4487C;
wire g1687C;
wire g2939C;
wire g6739C;
wire g7060C;
wire g1580C;
wire g5725C;
wire g11615C;
wire g2544C;
wire g11252C;
wire g5532C;
wire g3771C;
wire g11153C;
wire g9872C;
wire g9680C;
wire g9905C;
wire g7739C;
wire g6321C;
wire g8386C;
wire g8975C;
wire g2306C;
wire g6625C;
wire g7937C;
wire g8303C;
wire g8170C;
wire g5706C;
wire g2756C;
wire g8643C;
wire g8821C;
wire g5225C;
wire g10946C;
wire g4169C;
wire g5029C;
wire g11164C;
wire g4007C;
wire g1756C;
wire g4059C;
wire g1027C;
wire g4868C;
wire g5675C;
wire g4718C;
wire g10682C;
wire g6687C;
wire g682C;
wire g7704C;
wire g525C;
wire g1019C;
wire g4261C;
wire g3422C;
wire g5745C;
wire g8387C;
wire g7954C;
wire g11283C;
wire g8298C;
wire g8461C;
wire g10760C;
wire g11480C;
wire g6626C;
wire g6341C;
wire g10506C;
wire g16C;
wire g9648C;
wire g7453C;
wire g5995C;
wire g6645C;
wire g5707C;
wire g7548C;
wire g833C;
wire g11091C;
wire g496C;
wire g11174C;
wire g8403C;
wire g1250C;
wire g8605C;
wire g8841C;
wire g1914C;
wire g6879C;
wire g8763C;
wire g4502C;
wire g9702C;
wire g9839C;
wire g5841C;
wire g6358C;
wire g5575C;
wire g8107C;
wire g10240C;
wire g11192C;
wire g9618C;
wire g5539C;
wire g8416C;
wire g275C;
wire g9693C;
wire g11553C;
wire g7557C;
wire g1098C;
wire g5268C;
wire g9107C;
wire g10633C;
wire g7894C;
wire g8654C;
wire g9621C;
wire g5819C;
wire g6794C;
wire g3412C;
wire g7661C;
wire g2800C;
wire g3268C;
wire g9908C;
wire g3429C;
wire g351C;
wire g6628C;
wire g5470C;
wire g7526C;
wire g2204C;
wire g1482C;
wire g5025C;
wire g4921C;
wire g6204C;
wire g1750C;
wire g4048C;
wire g8935C;
wire g2525C;
wire g9593C;
wire g4827C;
wire g10701C;
wire g10733C;
wire g10777C;
wire g8130C;
wire g9955C;
wire g9965C;
wire g1710C;
wire g3684C;
wire g947C;
wire g11213C;
wire g1462C;
wire g5006C;
wire g9912C;
wire g9933C;
wire g8407C;
wire g8554C;
wire g9641C;
wire g6323C;
wire g10646C;
wire g10766C;
wire g6666C;
wire g4994C;
wire g5103C;
wire g3717C;
wire g11592C;
wire g1905C;
wire g6875C;
wire g9658C;
wire g6207C;
wire g6530C;
wire g8199C;
wire g7265C;
wire g9735C;
wire g9835C;
wire g6655C;
wire g3875C;
wire g7384C;
wire g7970C;
wire g1624C;
wire g5491C;
wire g8949C;
wire g11152C;
wire g9611C;
wire g2804C;
wire g6410C;
wire g10451C;
wire g4397C;
wire g5398C;
wire g7224C;
wire g5602C;
wire g6884C;
wire g8964C;
wire g11413C;
wire g1415C;
wire g4950C;
wire g5535C;
wire g6772C;
wire g7277C;
wire g8301C;
wire g8463C;
wire g2511C;
wire g10728C;
wire g6618C;
wire g6235C;
wire g6355C;
wire g3626C;
wire g4723C;
wire g8720C;
wire g6693C;
wire g11020C;
wire g1314C;
wire g11583C;
wire g8118C;
wire g8167C;
wire g7892C;
wire g8652C;
wire g5721C;
wire g10362C;
wire g10367C;
wire g9901C;
wire g290C;
wire g6792C;
wire g11282C;
wire g7945C;
wire g11302C;
wire g521C;
wire g3634C;
wire g11105C;
wire g8471C;
wire g8598C;
wire g7140C;
wire g9600C;
wire g1604C;
wire g9864C;
wire g11613C;
wire g5188C;
wire g7435C;
wire g7876C;
wire g1280C;
wire g4058C;
wire g5809C;
wire g6776C;
wire g630C;
wire g10301C;
wire g354C;
wire g4505C;
wire g17C;
wire g9623C;
wire g10739C;
wire g391C;
wire g11027C;
wire g10738C;
wire g8558C;
wire g8687C;
wire g6360C;
wire g1564C;
wire g9871C;
wire g5108C;
wire g11248C;
wire g4992C;
wire g11552C;
wire g944C;
wire g9651C;
wire g11204C;
wire g7824C;
wire g1133C;
wire g5115C;
wire g7102C;
wire g968C;
wire g9384C;
wire g2561C;
wire g9700C;
wire g9754C;
wire g9838C;
wire g10594C;
wire g10661C;
wire g11321C;
wire g8879C;
wire g7621C;
wire g8962C;
wire g2272C;
wire g10715C;
wire g8659C;
wire g950C;
wire g9643C;
wire g8957C;
wire g1669C;
wire g5538C;
wire g1744C;
wire g4000C;
wire g4126C;
wire g4088C;
wire g4400C;
wire I5886C;
wire I5887C;
wire g486C;
wire g6238C;
wire g10727C;
wire g8174C;
wire g305C;
wire g5067C;
wire g1512C;
wire g5418C;
wire g10297C;
wire g6353C;
wire g386C;
wire g11026C;
wire g11212C;
wire g4828C;
wire g6744C;
wire g1923C;
wire g10671C;
wire g2517C;
wire g4383C;
wire g4297C;
wire g5256C;
wire g4220C;
wire g8252C;
wire g8380C;
wire g7071C;
wire g9613C;
wire g8933C;
wire g5181C;
wire g7948C;
wire g324C;
wire g11149C;
wire g1601C;
wire g9862C;
wire g11387C;
wire g7955C;
wire g4161C;
wire g2321C;
wire g11148C;
wire g9712C;
wire g8931C;
wire g378C;
wire g11097C;
wire g3819C;
wire g2963C;
wire g11104C;
wire g1059C;
wire g6092C;
wire g4999C;
wire g4976C;
wire g632C;
wire g6858C;
wire g7409C;
wire g4103C;
wire I6309C;
wire g5944C;
wire g6580C;
wire g1056C;
wire g5631C;
wire g9414C;
wire g9660C;
wire g9926C;
wire g9946C;
wire I6331C;
wire g481C;
wire g9885C;
wire g9673C;
wire g9903C;
wire g10625C;
wire g6623C;
wire g11228C;
wire g11011C;
wire g1941C;
wire g6889C;
wire g7523C;
wire g7822C;
wire g8123C;
wire g11582C;
wire g4316C;
wire g3625C;
wire g10969C;
wire g5041C;
wire g9335C;
wire g9727C;
wire g9831C;
wire g9422C;
wire g4588C;
wire g8511C;
wire g8648C;
wire g8875C;
wire g5168C;
wire g7503C;
wire g7895C;
wire g8655C;
wire g1062C;
wire g4914C;
wire g9927C;
wire g9947C;
wire g1555C;
wire g5772C;
wire g1666C;
wire g5531C;
wire g5036C;
wire g10503C;
wire g7738C;
wire g8010C;
wire g8410C;
wire g5608C;
wire g6231C;
wire g10581C;
wire g10364C;
wire g10450C;
wire g2132C;
wire g2379C;
wire g9653C;
wire g1515C;
wire g10818C;
wire g8172C;
wire g10429C;
wire g5074C;
wire g1558C;
wire g9869C;
wire g10635C;
wire g10741C;
wire g8693C;
wire g5480C;
wire g3766C;
wire g4581C;
wire g2981C;
wire g8409C;
wire g8555C;
wire g9364C;
wire g506C;
wire g8994C;
wire g11299C;
wire g6592C;
wire g7958C;
wire g1474C;
wire g4995C;
wire g4079C;
wire g2264C;
wire g745C;
wire g2160C;
wire g3257C;
wire I6310C;
wire g1470C;
wire g5000C;
wire g3301C;
wire g1478C;
wire I5084C;
wire g1727C;
wire g9412C;
wire g1330C;
wire g9389C;
wire g10567C;
wire g10706C;
wire g10366C;
wire g10447C;
wire g10446C;
wire g10533C;
wire g5220C;
wire g10624C;
wire g10300C;
wire g5023C;
wire g4432C;
wire g4053C;
wire g7596C;
wire g1639C;
wire g5588C;
wire g6074C;
wire g9953C;
wire g9963C;
wire g3089C;
wire g3772C;
wire g5051C;
wire g8724C;
wire g4157C;
wire g1583C;
wire g9707C;
wire g8878C;
wire g10639C;
wire g10763C;
wire g6777C;
wire g8109C;
wire g7511C;
wire g7898C;
wire g11271C;
wire g11461C;
wire g5732C;
wire g315C;
wire g11145C;
wire g411C;
wire g11031C;
wire g1607C;
wire g9865C;
wire g1531C;
wire g9715C;
wire g9604C;
wire g8647C;
wire g8799C;
wire g11198C;
wire g6873C;
wire g6632C;
wire g6095C;
wire g9729C;
wire g9833C;
wire g1038C;
wire g6102C;
wire g7819C;
wire g11280C;
wire g7088C;
wire g9584C;
wire g9896C;
wire g8209C;
wire g6752C;
wire g11161C;
wire g8947C;
wire g5681C;
wire g7951C;
wire g9419C;
wire g1724C;
wire g5533C;
wire g8936C;
wire g178C;
wire g10670C;
wire g829C;
wire g11087C;
wire g4949C;
wire g5851C;
wire g6364C;
wire g7825C;
wire g1304C;
wire g10667C;
wire g7136C;
wire g339C;
wire g6532C;
wire g9385C;
wire g1436C;
wire g1440C;
wire g1448C;
wire g1137C;
wire g9897C;
wire g9425C;
wire g3383C;
wire g1035C;
wire g5601C;
wire g7943C;
wire g11171C;
wire I6631C;
wire g6064C;
wire g7230C;
wire g1648C;
wire g4952C;
wire g266C;
wire g6787C;
wire g8968C;
wire g10306C;
wire g11459C;
wire g538C;
wire g11458C;
wire g5739C;
wire g7496C;
wire g4986C;
wire g5187C;
wire g11010C;
wire g1741C;
wire g3999C;
wire g8175C;
wire g8722C;
wire g5590C;
wire g7471C;
wire g7891C;
wire g8651C;
wire g5479C;
wire g11599C;
wire g6684C;
wire g6745C;
wire g357C;
wire g6639C;
wire g3696C;
wire g4503C;
wire g6791C;
wire g8180C;
wire g1092C;
wire g4224C;
wire g5501C;
wire g8602C;
wire g8838C;
wire g10666C;
wire g309C;
wire g11158C;
wire g9602C;
wire g5704C;
wire g3879C;
wire g4617C;
wire g9868C;
wire g11295C;
wire g11144C;
wire g1540C;
wire g9718C;
wire g3434C;
wire g4987C;
wire g1270C;
wire g1065C;
wire g6098C;
wire g9582C;
wire g3533C;
wire g8104C;
wire g1733C;
wire g9415C;
wire g8377C;
wire g8499C;
wire g9664C;
wire g9413C;
wire g3584C;
wire g6162C;
wire g1508C;
wire g4991C;
wire g5846C;
wire g6362C;
wire g10685C;
wire g1153C;
wire g11023C;
wire g7598C;
wire g11224C;
wire g11571C;
wire g1520C;
wire g4959C;
wire g1633C;
wire g5626C;
wire g9920C;
wire g9940C;
wire g1086C;
wire g4876C;
wire g6730C;
wire g263C;
wire g9689C;
wire g10762C;
wire g1050C;
wire g6070C;
wire g9428C;
wire g1759C;
wire g9430C;
wire g8927C;
wire g7068C;
wire g7740C;
wire g8014C;
wire g11278C;
wire g5782C;
wire g4236C;
wire g11559C;
wire g9609C;
wire g11558C;
wire g6087C;
wire g10751C;
wire g10655C;
wire g10772C;
wire g8135C;
wire g11544C;
wire g5084C;
wire g8382C;
wire g10230C;
wire g7241C;
wire g3942C;
wire g10638C;
wire g4064C;
wire g1321C;
wire g9365C;
wire g9738C;
wire g9579C;
wire g9861C;
wire g11255C;
wire g11189C;
wire g10510C;
wire g2917C;
wire g11188C;
wire g9846C;
wire g1878C;
wire g7818C;
wire g11460C;
wire g11030C;
wire g841C;
wire g11093C;
wire g7478C;
wire g7893C;
wire g8653C;
wire g10442C;
wire g6535C;
wire g8102C;
wire g1490C;
wire g1494C;
wire I5085C;
wire g3912C;
wire g7186C;
wire g4489C;
wire g9662C;
wire g9418C;
wire g959C;
wire g11218C;
wire g1121C;
wire g10643C;
wire g10746C;
wire g7125C;
wire g7821C;
wire g6246C;
wire g8963C;
wire g7533C;
wire g10237C;
wire g7939C;
wire g8638C;
wire g8786C;
wire g10684C;
wire g11455C;
wire g8364C;
wire g2990C;
wire g9847C;
wire g7584C;
wire g5617C;
wire g5981C;
wire g5789C;
wire g4009C;
wire g11277C;
wire g6472C;
wire g6940C;
wire g6760C;
wire g7061C;
wire g11595C;
wire g5771C;
wire g8405C;
wire g8553C;
wire g4836C;
wire g5547C;
wire g4967C;
wire g342C;
wire g6671C;
wire g7200C;
wire g382C;
wire g7046C;
wire g999C;
wire g4229C;
wire g8389C;
wire g6430C;
wire g4993C;
wire g6247C;
wire g11170C;
wire g7145C;
wire g5738C;
wire g3998C;
wire g6741C;
wire g11167C;
wire g11194C;
wire g1333C;
wire g11589C;
wire g4431C;
wire g7536C;
wire g9585C;
wire g2957C;
wire g11588C;
wire g5690C;
wire g6883C;
wire g1068C;
wire g4837C;
wire g8641C;
wire g8791C;
wire g6217C;
wire g444C;
wire g11022C;
wire g4168C;
wire g5915C;
wire g511C;
wire g5110C;
wire g11254C;
wire g7567C;
wire g3273C;
wire g4392C;
wire g1592C;
wire g9856C;
wire g9411C;
wire g5002C;
wire g857C;
wire g11101C;
wire g11177C;
wire g11560C;
wire g8098C;
wire g3970C;
wire g4941C;
wire g366C;
wire g6662C;
wire g7935C;
wire g6067C;
wire g9740C;
wire g9863C;
wire g174C;
wire g170C;
wire g6758C;
wire g6994C;
wire g1589C;
wire g1007C;
wire g4252C;
wire g542C;
wire g11166C;
wire g7130C;
wire g5179C;
wire g11009C;
wire g7542C;
wire g5171C;
wire g11008C;
wire g1209C;
wire g3516C;
wire g7573C;
wire g3987C;
wire g491C;
wire g11555C;
wire g9734C;
wire g9569C;
wire g9857C;
wire g8728C;
wire g8730C;
wire g8185C;
wire g1610C;
wire g8385C;
wire g7902C;
wire g4073C;
wire g8070C;
wire g5731C;
wire g11238C;
wire g1125C;
wire g8308C;
wire g8470C;
wire g5489C;
wire g3991C;
wire g166C;
wire g7823C;
wire g4069C;
wire g1317C;
wire g11176C;
wire g837C;
wire g11092C;
wire g330C;
wire g11154C;
wire g7C;
wire g9608C;
wire g11637C;
wire g2091C;
wire g8406C;
wire g5254C;
wire g8612C;
wire g9588C;
wire g8742C;
wire g8801C;
wire g7063C;
wire g10303C;
wire g1486C;
wire g5009C;
wire g9665C;
wire g8748C;
wire g11215C;
wire g10750C;
wire g3818C;
wire g5769C;
wire g6673C;
wire g1255C;
wire g7720C;
wire g4609C;
wire g7547C;
wire g7971C;
wire g11288C;
wire g7599C;
wire g6058C;
wire g4106C;
wire g6743C;
wire g6890C;
wire g7269C;
wire g7549C;
wire g8169C;
wire g11304C;
wire g9924C;
wire g9944C;
wire g7592C;
wire g8718C;
wire g8616C;
wire g9316C;
wire g7625C;
wire g8644C;
wire g8793C;
wire g2940C;
wire g11624C;
wire g2947C;
wire g10949C;
wire g3563C;
wire g2223C;
wire g10948C;
wire g7846C;
wire g8246C;
wire g5788C;
wire g4008C;
wire g9596C;
wire g5249C;
wire g11585C;
wire g4972C;
wire g11554C;
wire g7096C;
wire g10673C;
wire g2493C;
wire g4806C;
wire g9915C;
wire g9936C;
wire g1660C;
wire g2910C;
wire g9317C;
wire g10853C;
wire g10933C;
wire g8177C;
wire g8388C;
wire g1117C;
wire g7141C;
wire g10508C;
wire g4230C;
wire g10634C;
wire g9192C;
wire g9601C;
wire g6326C;
wire g700C;
wire g7710C;
wire g7375C;
wire g8028C;
wire g5640C;
wire g5031C;
wire g4550C;
wire g7879C;
wire g7962C;
wire g9597C;
wire g631C;
wire g5005C;
wire g6423C;
wire g8108C;
wire g3322C;
wire g5911C;
wire g9916C;
wire g9937C;
wire g9704C;
wire g9747C;
wire g9840C;
wire g10723C;
wire g8217C;
wire g5209C;
wire g11013C;
wire g9390C;
wire g11214C;
wire g6327C;
wire g1149C;
wire g5796C;
wire g5473C;
wire g5038C;
wire g6346C;
wire g6633C;
wire g5119C;
wire g11005C;
wire g8365C;
wire g7558C;
wire g4481C;
wire g4097C;
wire g7588C;
wire g4497C;
wire g9922C;
wire g9942C;
wire g6696C;
wire g5118C;
wire g1850C;
wire g10665C;
wire g10731C;
wire g8552C;
wire g8827C;
wire g5540C;
wire g1403C;
wire g4960C;
wire g8615C;
wire g8846C;
wire g5983C;
wire g182C;
wire g6240C;
wire g7931C;
wire g853C;
wire g11100C;
wire g11235C;
wire g5199C;
wire g6316C;
wire g7515C;
wire g5781C;
wire g7742C;
wire g8018C;
wire g2950C;
wire g5510C;
wire g6347C;
wire g962C;
wire g9357C;
wire g11407C;
wire g10743C;
wire g5259C;
wire g5694C;
wire g10769C;
wire g11584C;
wire g4932C;
wire g10649C;
wire g10768C;
wire g4068C;
wire g6317C;
wire g4276C;
wire g5215C;
wire g6775C;
wire g10662C;
wire g8101C;
wire g3204C;
wire g5318C;
wire g5825C;
wire g7457C;
wire g7884C;
wire g1292C;
wire g3974C;
wire g9929C;
wire g9949C;
wire g10778C;
wire g7524C;
wire g6079C;
wire g7235C;
wire g9603C;
wire g9726C;
wire g9850C;
wire g7988C;
wire g5228C;
wire g5587C;
wire g5934C;
wire g8168C;
wire g9583C;
wire g10672C;
wire g8627C;
wire g635C;
wire g8309C;
wire g10449C;
wire g11273C;
wire g8734C;
wire g5913C;
wire g4572C;
wire g6363C;
wire g11463C;
wire g718C;
wire g8074C;
wire g1166C;
wire g8383C;
wire g8474C;
wire g11234C;
wire g4483C;
wire g11491C;
wire g5097C;
wire g5726C;
wire g5497C;
wire g7933C;
wire g9C;
wire g9617C;
wire g9873C;
wire g9906C;
wire g5196C;
wire g11012C;
wire g7050C;
wire g10849C;
wire g10971C;
wire g8400C;
wire g1169C;
wire g4345C;
wire g9925C;
wire g9945C;
wire g5028C;
wire g7271C;
wire g9709C;
wire g1003C;
wire g4223C;
wire g10497C;
wire g10716C;
wire g11247C;
wire g6661C;
wire g11173C;
wire g6075C;
wire g7367C;
wire g8023C;
wire g9888C;
wire g9907C;
wire g10582C;
wire g5746C;
wire g9950C;
wire g9959C;
wire g7674C;
wire g9690C;
wire g5703C;
wire g360C;
wire g4522C;
wire g4115C;
wire g7075C;
wire g10627C;
wire g4047C;
wire g2944C;
wire g6646C;
wire g7132C;
wire g11029C;
wire g7572C;
wire g8127C;
wire g7209C;
wire g11028C;
wire g10742C;
wire g8880C;
wire g10681C;
wire g9663C;
wire g5349C;
wire g8732C;
wire g3807C;
wire g3860C;
wire g5848C;
wire g8411C;
wire g8508C;
wire g8072C;
wire g5699C;
wire g11240C;
wire g6105C;
wire g6616C;
wire g10690C;
wire g7582C;
wire g9590C;
wire g4128C;
wire g6404C;
wire g6647C;
wire g10504C;
wire g9657C;
wire g4542C;
wire g1163C;
wire g5524C;
wire g9899C;
wire g7736C;
wire g10626C;
wire g6320C;
wire g7623C;
wire g10299C;
wire g7889C;
wire g10298C;
wire g8413C;
wire g3979C;
wire g1848C;
wire g5211C;
wire g4512C;
wire g7722C;
wire g9714C;
wire g9522C;
wire g9844C;
wire g1141C;
wire g5993C;
wire g5026C;
wire g8705C;
wire g10737C;
wire g10232C;
wire g6771C;
wire g5170C;
wire g8117C;
wire g9956C;
wire g9966C;
wire g5280C;
wire g7139C;
wire g11099C;
wire g6892C;
wire g9705C;
wire g10512C;
wire g849C;
wire g11098C;
wire g8628C;
wire g5544C;
wire g11272C;
wire g1621C;
wire g5483C;
wire g9928C;
wire g9948C;
wire g4063C;
wire g11462C;
wire g6738C;
wire g7593C;
wire g11032C;
wire g10445C;
wire g8882C;
wire g10316C;
wire g5756C;
wire g1023C;
wire g4720C;
wire g9409C;
wire g8929C;
wire g6876C;
wire g4989C;
wire g9737C;
wire g9836C;
wire g6061C;
wire g8268C;
wire g6465C;
wire g1466C;
wire g5003C;
wire g9957C;
wire g9967C;
wire g5145C;
wire g4971C;
wire g10753C;
wire g5695C;
wire g7613C;
wire g10736C;
wire g11220C;
wire g7444C;
wire g4670C;
wire g4253C;
wire g7960C;
wire g8163C;
wire g10764C;
wire g5757C;
wire g7385C;
wire g8032C;
wire g2988C;
wire g11591C;
wire g7583C;
wire g321C;
wire g11147C;
wire g5522C;
wire g1394C;
wire g9697C;
wire g9751C;
wire g9837C;
wire g9620C;
wire g327C;
wire g11151C;
wire g11172C;
wire g7885C;
wire g5595C;
wire g5537C;
wire g9708C;
wire g9516C;
wire g9842C;
wire g4141C;
wire g4341C;
wire g7679C;
wire g7378C;
wire g5612C;
wire g7135C;
wire g10970C;
wire g11025C;
wire g9730C;
wire g9854C;
wire g7182C;
wire g9921C;
wire g9941C;
wire g6194C;
wire g1651C;
wire g4962C;
wire g4358C;
wire g4803C;
wire g8549C;
wire g8683C;
wire g1113C;
wire g5224C;
wire g8778C;
wire g11281C;
wire g318C;
wire g11146C;
wire g2948C;
wire g3904C;
wire g8075C;
wire g9723C;
wire g9829C;
wire g7184C;
wire g11246C;
wire g5837C;
wire g6350C;
wire g2555C;
wire g5902C;
wire g1765C;
wire g6438C;
wire g5512C;
wire g5090C;
wire g7719C;
wire g3695C;
wire g7587C;
wire g9610C;
wire g3536C;
wire g8881C;
wire g4559C;
wire g10549C;
wire g10561C;
wire g5698C;
wire g11226C;
wire g10295C;
wire g5260C;
wire g10680C;
wire g1853C;
wire g11538C;
wire g11551C;
wire g9849C;
wire g5279C;
wire g8404C;
wire g5720C;
wire g11318C;
wire g11297C;
wire g9898C;
wire g9510C;
wire g7297C;
wire g7963C;
wire g9759C;
wire g9803C;
wire g11338C;
wire g8435C;
wire g6124C;
wire I5600C;
wire g11257C;
wire g11256C;
wire g3107C;
wire g2167C;
wire I14866C;
wire g4997C;
wire g10291C;
wire g6122C;
wire g9509C;
wire g5227C;
wire I15054C;
wire g11269C;
wire g5555C;
wire g11268C;
wire g11335C;
wire g8249C;
wire g9882C;
wire I15210C;
wire g2102C;
wire g2099C;
wire g2096C;
wire g2088C;
wire I5805C;
wire g11443C;
wire g8431C;
wire g8286C;
wire g7290C;
wire g8287C;
wire g7301C;
wire g8259C;
wire g11334C;
wire g10805C;
wire I15214C;
wire I15215C;
wire g11265C;
wire g8322C;
wire g8433C;
wire g8248C;
wire g8154C;
wire g2405C;
wire g2389C;
wire g2380C;
wire g2372C;
wire I6351C;
wire I16427C;
wire g7303C;
wire g2862C;
wire g2515C;
wire g4052C;
wire I14858C;
wire g11264C;
wire I15209C;
wire g1570C;
wire g2528C;
wire g2522C;
wire g9515C;
wire g7294C;
wire g3118C;
wire g2180C;
wire I5571C;
wire I5599C;
wire g2514C;
wire g11327C;
wire I5629C;
wire I5363C;
wire g2315C;
wire g8159C;
wire g11326C;
wire I16148C;
wire I16149C;
wire g10521C;
wire g7292C;
wire g8417C;
wire I14855C;
wire g9878C;
wire I15205C;
wire I15051C;
wire g8823C;
wire g8148C;
wire g2863C;
wire g2516C;
wire g7299C;
wire g9511C;
wire g9654C;
wire I15224C;
wire I15225C;
wire g8253C;
wire I15171C;
wire I15172C;
wire I15204C;
wire g10472C;
wire g10470C;
wire g10468C;
wire g10467C;
wire g10386C;
wire g10384C;
wire g10476C;
wire g10474C;
wire g8158C;
wire g11331C;
wire g7295C;
wire g8284C;
wire g1393C;
wire I5357C;
wire g9758C;
wire I5626C;
wire g7298C;
wire g8282C;
wire I15057C;
wire I15219C;
wire I15220C;
wire I14862C;
wire g2521C;
wire g9591C;
wire g9757C;
wire g11261C;
wire g9815C;
wire I14835C;
wire g126C;
wire g10479C;
wire g10478C;
wire g10477C;
wire g10475C;
wire I16161C;
wire g2353C;
wire I5804C;
wire g7291C;
wire I15199C;
wire g11330C;
wire g8153C;
wire g9881C;
wire g11259C;
wire g11258C;
wire g9426C;
wire g9423C;
wire g11337C;
wire g8262C;
wire g8285C;
wire I5570C;
wire g2499C;
wire g11336C;
wire g7293C;
wire g9388C;
wire g11260C;
wire g10807C;
wire g8288C;
wire g10394C;
wire g10392C;
wire g10482C;
wire g10481C;
wire I16160C;
wire g9589C;
wire g11270C;
wire g11267C;
wire g1959C;
wire g9667C;
wire I14827C;
wire g9391C;
wire I5358C;
wire g2309C;
wire g11266C;
wire g8429C;
wire g8281C;
wire g9876C;
wire I15177C;
wire g5186C;
wire I6350C;
wire g1527C;
wire g8162C;
wire I14779C;
wire I5351C;
wire I5352C;
wire g2305C;
wire I15176C;
wire g9879C;
wire g8283C;
wire g11333C;
wire g10562C;
wire g9606C;
wire I14822C;
wire g9880C;
wire I15200C;
wire g8428C;
wire g8430C;
wire g8247C;
wire I5576C;
wire g4476C;
wire I5649C;
wire g2538C;
wire g11329C;
wire g11328C;
wire g9605C;
wire g9363C;
wire g7300C;
wire I14831C;
wire g8263C;
wire g11263C;
wire g5780C;
wire g11332C;
wire I15048C;
wire g9647C;
wire I14602C;
wire I15033C;
wire g2445C;
wire g2437C;
wire g2433C;
wire g2419C;
wire g11325C;
wire I5366C;
wire g9506C;
wire g8161C;
wire g2316C;
wire g4675C;
wire g8434C;
wire g11262C;
wire g9387C;
wire I15045C;
wire g11324C;
wire g2501C;
wire g9877C;
wire g10529C;
wire g8432C;
wire g9874C;
wire g8157C;
wire g6899C;
wire g9646C;
wire g7302C;
wire g2111C;
wire g2109C;
wire g2106C;
wire g2104C;
wire g7296C;
wire I5612C;
wire I5613C;
wire I5591C;
wire I5593C;
wire g8839C;
wire g8970C;
wire I10519C;
wire I11278C;
wire I11279C;
wire g3978C;
wire I5263C;
wire I5264C;
wire g4278C;
wire I8640C;
wire g2943C;
wire I6760C;
wire I6761C;
wire g11418C;
wire g11416C;
wire I17400C;
wire I5449C;
wire I5450C;
wire I16058C;
wire I16060C;
wire g2938C;
wire I6746C;
wire I11973C;
wire I11975C;
wire I12136C;
wire I11935C;
wire I11937C;
wire I6167C;
wire I6168C;
wire g2959C;
wire g2120C;
wire g2115C;
wire I5878C;
wire I5619C;
wire I5620C;
wire g5552C;
wire I6467C;
wire I6468C;
wire g4672C;
wire I8795C;
wire I8796C;
wire I15891C;
wire I15892C;
wire I5611C;
wire g8738C;
wire I6714C;
wire I6716C;
wire g3460C;
wire I7683C;
wire I7685C;
wire I12106C;
wire I12108C;
wire I6747C;
wire I5230C;
wire I5231C;
wire g2236C;
wire I12075C;
wire I12076C;
wire I15870C;
wire I16065C;
wire I16067C;
wire I7562C;
wire I13529C;
wire I13531C;
wire I8797C;
wire I17584C;
wire I11936C;
wire I15256C;
wire I15257C;
wire I13505C;
wire I13506C;
wire g8502C;
wire g8501C;
wire g8824C;
wire I6186C;
wire I17504C;
wire I17505C;
wire g11496C;
wire I15999C;
wire I16001C;
wire g2215C;
wire I6124C;
wire I6125C;
wire I11907C;
wire I11909C;
wire I12038C;
wire I12040C;
wire I13907C;
wire I13909C;
wire I6771C;
wire I6772C;
wire I11908C;
wire I16008C;
wire I16009C;
wire I13908C;
wire I7034C;
wire I7035C;
wire I8650C;
wire I9947C;
wire I9948C;
wire g10428C;
wire I16066C;
wire I6144C;
wire I6145C;
wire I11241C;
wire I11242C;
wire I15993C;
wire I15994C;
wire I6187C;
wire g6027C;
wire I5500C;
wire I11974C;
wire I12060C;
wire I12062C;
wire I8771C;
wire I8772C;
wire I5184C;
wire I13293C;
wire I6199C;
wire I6200C;
wire I13265C;
wire I5023C;
wire I5024C;
wire I7863C;
wire I13991C;
wire I13992C;
wire I13660C;
wire I13661C;
wire I6143C;
wire I13990C;
wire I11508C;
wire I11510C;
wire g5034C;
wire I5229C;
wire I12045C;
wire I12047C;
wire I10769C;
wire I10771C;
wire I16045C;
wire I16046C;
wire I12061C;
wire I5104C;
wire I13530C;
wire I6447C;
wire I4954C;
wire I4956C;
wire g3530C;
wire I8479C;
wire I8481C;
wire I8739C;
wire I8740C;
wire I6879C;
wire I6880C;
wire I15430C;
wire I15431C;
wire I12019C;
wire I12020C;
wire I16331C;
wire I16332C;
wire I16467C;
wire I16469C;
wire I5013C;
wire I5014C;
wire I13521C;
wire I13523C;
wire I16037C;
wire I16039C;
wire I16468C;
wire I12046C;
wire I16038C;
wire g4374C;
wire I8676C;
wire I12113C;
wire g4616C;
wire I8761C;
wire I15992C;
wire I5034C;
wire I5036C;
wire g8843C;
wire I14263C;
wire I13249C;
wire I13250C;
wire I5135C;
wire I5485C;
wire I5486C;
wire I7033C;
wire I15441C;
wire I15443C;
wire I6166C;
wire g4267C;
wire I8624C;
wire I16015C;
wire I8677C;
wire g4234C;
wire I8575C;
wire I8576C;
wire g9204C;
wire I14612C;
wire I14613C;
wire g4601C;
wire I8715C;
wire I8716C;
wire I6715C;
wire I13514C;
wire I13515C;
wire I12002C;
wire I12003C;
wire I5127C;
wire I5128C;
wire g2177C;
wire I8577C;
wire g11414C;
wire I17393C;
wire I17395C;
wire I11280C;
wire I5265C;
wire I6988C;
wire I6989C;
wire I13272C;
wire I13274C;
wire I10507C;
wire I5164C;
wire I14443C;
wire I14444C;
wire I9557C;
wire I9559C;
wire I5592C;
wire I13077C;
wire I13078C;
wire I8717C;
wire I5295C;
wire I5296C;
wire I8625C;
wire I8626C;
wire I4911C;
wire I4912C;
wire I16000C;
wire I5371C;
wire I5185C;
wire I5186C;
wire I5675C;
wire g4218C;
wire I8543C;
wire I8544C;
wire I10520C;
wire I10521C;
wire I5297C;
wire I13537C;
wire I13283C;
wire g4749C;
wire I11980C;
wire I11982C;
wire g4873C;
wire I8513C;
wire I8514C;
wire I13089C;
wire I13091C;
wire I6126C;
wire g10302C;
wire I15906C;
wire I15908C;
wire I8763C;
wire g8506C;
wire g8825C;
wire I16007C;
wire g2107C;
wire g2105C;
wire I5865C;
wire I5604C;
wire I5517C;
wire I5518C;
wire I6109C;
wire I6111C;
wire I4929C;
wire I4930C;
wire I13522C;
wire I10770C;
wire I5538C;
wire I5539C;
wire g11415C;
wire I17394C;
wire I13552C;
wire I13553C;
wire I8642C;
wire I17296C;
wire I17297C;
wire I14278C;
wire I14279C;
wire I4910C;
wire I6792C;
wire I6794C;
wire I5484C;
wire I15442C;
wire I10931C;
wire I10932C;
wire I8779C;
wire I8780C;
wire g2354C;
wire g10043C;
wire g10153C;
wire I15615C;
wire I17281C;
wire I5468C;
wire I5470C;
wire I11509C;
wire I5025C;
wire I14270C;
wire I14272C;
wire I6208C;
wire I6209C;
wire I17288C;
wire I17290C;
wire I7563C;
wire I7564C;
wire I5005C;
wire I5006C;
wire I12126C;
wire I12128C;
wire I5105C;
wire I6322C;
wire I6323C;
wire I12093C;
wire I12094C;
wire g2776C;
wire I6664C;
wire I6666C;
wire I6762C;
wire g3623C;
wire I5373C;
wire I8527C;
wire I8529C;
wire I5282C;
wire I5283C;
wire I7223C;
wire I7224C;
wire I5007C;
wire I5459C;
wire I17295C;
wire I5015C;
wire I14264C;
wire I14265C;
wire I16072C;
wire I16073C;
wire g3205C;
wire I8652C;
wire I9558C;
wire I5202C;
wire I5203C;
wire I6806C;
wire I6807C;
wire I6469C;
wire I12143C;
wire I12145C;
wire I12127C;
wire I13300C;
wire I13302C;
wire I5502C;
wire I9574C;
wire I6448C;
wire I6449C;
wire I8669C;
wire I8670C;
wire I15451C;
wire I15453C;
wire I7875C;
wire I7876C;
wire I14202C;
wire I14203C;
wire g10149C;
wire g10144C;
wire I15607C;
wire I5324C;
wire I5325C;
wire I8738C;
wire g10434C;
wire g5859C;
wire I8604C;
wire I8606C;
wire I12085C;
wire I12087C;
wire I13248C;
wire I4979C;
wire I4980C;
wire I12067C;
wire I12069C;
wire g8942C;
wire I12068C;
wire I17503C;
wire I7877C;
wire I5165C;
wire I6287C;
wire I6289C;
wire I6777C;
wire I8562C;
wire I8563C;
wire I15890C;
wire g8006C;
wire I13090C;
wire I17460C;
wire I17461C;
wire g11474C;
wire I13513C;
wire I4986C;
wire I4987C;
wire I5204C;
wire I13504C;
wire I6207C;
wire I12086C;
wire I8545C;
wire I8178C;
wire I8180C;
wire I8589C;
wire I8591C;
wire I10930C;
wire I17402C;
wire I13294C;
wire I13295C;
wire I12144C;
wire g8757C;
wire g2961C;
wire I14209C;
wire I14211C;
wire I8515C;
wire I5316C;
wire I5317C;
wire I9946C;
wire g4613C;
wire I8750C;
wire I5605C;
wire I14204C;
wire I16051C;
wire g10360C;
wire g6037C;
wire I13858C;
wire I13859C;
wire I15872C;
wire g4879C;
wire I8528C;
wire I13901C;
wire I13902C;
wire g8542C;
wire I6836C;
wire I6838C;
wire I17305C;
wire I17307C;
wire g4538C;
wire I15452C;
wire I13857C;
wire I13765C;
wire I8671C;
wire I16044C;
wire g10363C;
wire g5360C;
wire I5106C;
wire g4677C;
wire I8803C;
wire I8804C;
wire I16016C;
wire I16017C;
wire I17485C;
wire I17487C;
wire I4995C;
wire I12092C;
wire I8678C;
wire I5126C;
wire I5372C;
wire I17306C;
wire I11995C;
wire I7225C;
wire I11261C;
wire g8545C;
wire I6110C;
wire I4941C;
wire I4942C;
wire I15899C;
wire I15900C;
wire g5527C;
wire g5350C;
wire I16079C;
wire I16081C;
wire I8641C;
wire I6176C;
wire I6178C;
wire I12074C;
wire I5451C;
wire I7322C;
wire I7323C;
wire I6288C;
wire I8179C;
wire I6805C;
wire I17486C;
wire I4928C;
wire I16330C;
wire I9575C;
wire I13886C;
wire I13887C;
wire I8787C;
wire I8788C;
wire I5315C;
wire g10285C;
wire I13867C;
wire I13869C;
wire I13868C;
wire I13258C;
wire I13259C;
wire g3261C;
wire I16074C;
wire I5136C;
wire I5137C;
wire I5460C;
wire I5461C;
wire I8605C;
wire I6770C;
wire I17401C;
wire g11449C;
wire g11448C;
wire g10231C;
wire I15716C;
wire I15717C;
wire I14210C;
wire I17567C;
wire I17569C;
wire I13876C;
wire I13878C;
wire I5606C;
wire I14442C;
wire I11996C;
wire I11997C;
wire I14277C;
wire I17568C;
wire I7321C;
wire I6990C;
wire g8847C;
wire I9006C;
wire I4985C;
wire I8651C;
wire I13544C;
wire I13545C;
wire I13894C;
wire I13895C;
wire I6136C;
wire I6138C;
wire I13076C;
wire g2205C;
wire I13260C;
wire I5501C;
wire I17586C;
wire I13900C;
wire I6201C;
wire g8826C;
wire I14216C;
wire I14217C;
wire I9007C;
wire I13559C;
wire I13561C;
wire g10229C;
wire I17492C;
wire I17493C;
wire I12214C;
wire I12215C;
wire I11262C;
wire I11263C;
wire I6225C;
wire I6226C;
wire I13307C;
wire I13309C;
wire I5676C;
wire I5677C;
wire I6826C;
wire I6827C;
wire g8190C;
wire I13308C;
wire I5879C;
wire I5880C;
wire g2792C;
wire g3061C;
wire I17585C;
wire I6881C;
wire I12138C;
wire g4605C;
wire I8728C;
wire I8729C;
wire I15871C;
wire I5866C;
wire I5867C;
wire I6793C;
wire I6487C;
wire I16080C;
wire I13893C;
wire I12115C;
wire I6748C;
wire I6224C;
wire I8805C;
wire I15878C;
wire I15880C;
wire I16030C;
wire I16031C;
wire I14271C;
wire I13267C;
wire I15616C;
wire I15617C;
wire I4964C;
wire I4966C;
wire I8752C;
wire I15432C;
wire g10438C;
wire g6032C;
wire g3011C;
wire I8480C;
wire I16086C;
wire I16087C;
wire g3734C;
wire I14218C;
wire I4955C;
wire g4639C;
wire I8786C;
wire g10480C;
wire I11914C;
wire I11915C;
wire g4619C;
wire I8770C;
wire I5516C;
wire g8541C;
wire I6188C;
wire I5891C;
wire I5892C;
wire I13766C;
wire I13767C;
wire I15258C;
wire I13266C;
wire I6825C;
wire I17283C;
wire g5277C;
wire I5035C;
wire g10359C;
wire I15879C;
wire I12114C;
wire I12107C;
wire g2500C;
wire g10430C;
wire g5999C;
wire I13285C;
wire I13877C;
wire I5893C;
wire g2795C;
wire I13560C;
wire g4259C;
wire I5166C;
wire I14614C;
wire I4965C;
wire I4943C;
wire I16023C;
wire I16059C;
wire g8737C;
wire I9576C;
wire I16052C;
wire I16053C;
wire I12004C;
wire g5573C;
wire I6837C;
wire I8730C;
wire I4978C;
wire I6177C;
wire I17051C;
wire I7864C;
wire I7865C;
wire I6665C;
wire I12216C;
wire I13554C;
wire I13284C;
wire I6137C;
wire I5529C;
wire I5530C;
wire I17282C;
wire I5618C;
wire I8662C;
wire I8664C;
wire I11916C;
wire g7717C;
wire I4971C;
wire I4972C;
wire I13273C;
wire I10509C;
wire I10508C;
wire I6778C;
wire I6779C;
wire I5469C;
wire g4251C;
wire I13546C;
wire I4996C;
wire I4997C;
wire I13539C;
wire I16032C;
wire I5323C;
wire I13538C;
wire I5540C;
wire I8778C;
wire g4286C;
wire I17052C;
wire I17053C;
wire I15898C;
wire g7978C;
wire g4227C;
wire I8561C;
wire I8762C;
wire I8751C;
wire I15907C;
wire I4973C;
wire I16024C;
wire I16025C;
wire g4455C;
wire I5341C;
wire I5342C;
wire I12137C;
wire I16088C;
wire g10483C;
wire I17289C;
wire g4630C;
wire I15609C;
wire I15608C;
wire g10436C;
wire g6023C;
wire I17459C;
wire I13301C;
wire I11981C;
wire I8663C;
wire I15718C;
wire I5284C;
wire g4607C;
wire g8840C;
wire g10441C;
wire g5345C;
wire g10432C;
wire g5938C;
wire I12021C;
wire I6489C;
wire I5528C;
wire I13659C;
wire I5343C;
wire I12039C;
wire I9008C;
wire I6488C;
wire I13888C;
wire I17494C;
wire I7684C;
wire g3221C;
wire I6324C;
wire I8590C;
wire I11243C;
wire g1737C;
wire g10324C;
wire g10239C;
wire g4974C;
wire g10322C;
wire g1736C;
wire g1955C;
wire g1956C;
wire g113C;
wire g1360C;
wire g1217C;
wire g755C;
wire g875C;
wire g1356C;
wire g874C;

assign test_soA= g73A;
assign test_soB= g73B;
assign test_soC= g73C;

INV_X1 FE_OFC370_g4525A (.ZN(FE_OFN370_g4525A),.A(FE_OFN368_g4525A));
INV_X1 FE_OFC369_g4525A (.ZN(FE_OFN369_g4525A),.A(FE_OFN368_g4525A));
INV_X1 FE_OFC368_g4525A (.ZN(FE_OFN368_g4525A),.A(FE_OFN362_g4525A));
BUF_X3 FE_OFC367_g3521A (.Z(FE_OFN367_g3521A),.A(FE_OFN366_g3521A));
BUF_X3 FE_OFC366_g3521A (.Z(FE_OFN366_g3521A),.A(FE_OFN358_g3521A));
BUF_X3 FE_OFC365_g5361A (.Z(FE_OFN365_g5361A),.A(FE_OFN356_g5361A));
BUF_X3 FE_OFC364_g3015A (.Z(FE_OFN364_g3015A),.A(FE_OFN348_g3015A));
BUF_X3 FE_OFC363_I5565A (.Z(FE_OFN363_I5565A),.A(FE_OFN343_I5565A));
INV_X1 FE_OFC362_g4525A (.ZN(FE_OFN362_g4525A),.A(FE_OFN360_g4525A));
INV_X1 FE_OFC360_g4525A (.ZN(FE_OFN360_g4525A),.A(FE_OFN339_g4525A));
BUF_X3 FE_OFC359_g18A (.Z(FE_OFN359_g18A),.A(FE_OFN324_g18A));
BUF_X3 FE_OFC358_g3521A (.Z(FE_OFN358_g3521A),.A(g3521A));
BUF_X3 FE_OFC357_g3521A (.Z(FE_OFN357_g3521A),.A(FE_OFN366_g3521A));
INV_X1 FE_OFC356_g5361A (.ZN(FE_OFN356_g5361A),.A(FE_OFN354_g5361A));
INV_X1 FE_OFC354_g5361A (.ZN(FE_OFN354_g5361A),.A(FE_OFN318_g5361A));
BUF_X3 FE_OFC353_g5117A (.Z(FE_OFN353_g5117A),.A(FE_OFN315_g5117A));
BUF_X3 FE_OFC352_g109A (.Z(FE_OFN352_g109A),.A(FE_OFN269_g109A));
BUF_X3 FE_OFC351_g3913A (.Z(FE_OFN351_g3913A),.A(FE_OFN302_g3913A));
BUF_X3 FE_OFC350_g3121A (.Z(FE_OFN350_g3121A),.A(FE_OFN155_g3121A));
BUF_X3 FE_OFC349_I6424A (.Z(FE_OFN349_I6424A),.A(FE_OFN308_I6424A));
BUF_X3 FE_OFC348_g3015A (.Z(FE_OFN348_g3015A),.A(FE_OFN298_g3015A));
BUF_X3 FE_OFC347_g3914A (.Z(FE_OFN347_g3914A),.A(FE_OFN296_g3914A));
BUF_X3 FE_OFC346_g4381A (.Z(FE_OFN346_g4381A),.A(g4381A));
BUF_X3 FE_OFC345_g3015A (.Z(FE_OFN345_g3015A),.A(FE_OFN297_g3015A));
BUF_X3 FE_OFC344_g3586A (.Z(FE_OFN344_g3586A),.A(FE_OFN287_g3586A));
INV_X1 FE_OFC343_I5565A (.ZN(FE_OFN343_I5565A),.A(FE_OFN340_I5565A));
INV_X1 FE_OFC340_I5565A (.ZN(FE_OFN340_I5565A),.A(FE_OFN233_I5565A));
INV_X1 FE_OFC339_g4525A (.ZN(FE_OFN339_g4525A),.A(FE_OFN337_g4525A));
INV_X1 FE_OFC337_g4525A (.ZN(FE_OFN337_g4525A),.A(g4525A));
BUF_X3 FE_OFC336_g1690A (.Z(FE_OFN336_g1690A),.A(FE_OFN245_g1690A));
BUF_X3 FE_OFC335_g4737A (.Z(FE_OFN335_g4737A),.A(g4737A));
BUF_X3 FE_OFC334_g7045A (.Z(FE_OFN334_g7045A),.A(g7045A));
BUF_X3 FE_OFC333_g4294A (.Z(FE_OFN333_g4294A),.A(g4294A));
BUF_X3 FE_OFC332_g8748A (.Z(FE_OFN332_g8748A),.A(g8748A));
BUF_X3 FE_OFC331_g8696A (.Z(FE_OFN331_g8696A),.A(g8696A));
BUF_X3 FE_OFC330_g7638A (.Z(FE_OFN330_g7638A),.A(FE_OFN189_g7638A));
BUF_X3 FE_OFC329_g8763A (.Z(FE_OFN329_g8763A),.A(g8763A));
BUF_X3 FE_OFC328_g8709A (.Z(FE_OFN328_g8709A),.A(g8709A));
BUF_X3 FE_OFC325_g18A (.Z(FE_OFN325_g18A),.A(FE_OFN359_g18A));
BUF_X3 FE_OFC324_g18A (.Z(FE_OFN324_g18A),.A(FE_OFN260_g18A));
BUF_X3 FE_OFC322_g4449A (.Z(FE_OFN322_g4449A),.A(g4449A));
BUF_X3 FE_OFC321_g5261A (.Z(FE_OFN321_g5261A),.A(g5261A));
BUF_X3 FE_OFC320_g5361A (.Z(FE_OFN320_g5361A),.A(FE_OFN319_g5361A));
BUF_X3 FE_OFC319_g5361A (.Z(FE_OFN319_g5361A),.A(FE_OFN166_g5361A));
INV_X1 FE_OFC318_g5361A (.ZN(FE_OFN318_g5361A),.A(FE_OFN316_g5361A));
INV_X1 FE_OFC316_g5361A (.ZN(FE_OFN316_g5361A),.A(FE_OFN168_g5361A));
INV_X1 FE_OFC315_g5117A (.ZN(FE_OFN315_g5117A),.A(FE_OFN312_g5117A));
INV_X1 FE_OFC312_g5117A (.ZN(FE_OFN312_g5117A),.A(g5117A));
BUF_X3 FE_OFC310_g4336A (.Z(FE_OFN310_g4336A),.A(g4336A));
BUF_X3 FE_OFC308_I6424A (.Z(FE_OFN308_I6424A),.A(FE_OFN160_I6424A));
BUF_X3 FE_OFC307_g4010A (.Z(FE_OFN307_g4010A),.A(g4010A));
BUF_X3 FE_OFC306_g5128A (.Z(FE_OFN306_g5128A),.A(g5128A));
BUF_X3 FE_OFC305_g5151A (.Z(FE_OFN305_g5151A),.A(FE_OFN304_g5151A));
BUF_X3 FE_OFC304_g5151A (.Z(FE_OFN304_g5151A),.A(FE_OFN176_g5151A));
BUF_X3 FE_OFC303_g4678A (.Z(FE_OFN303_g4678A),.A(g4678A));
BUF_X3 FE_OFC302_g3913A (.Z(FE_OFN302_g3913A),.A(g3913A));
BUF_X3 FE_OFC300_g4002A (.Z(FE_OFN300_g4002A),.A(g4002A));
BUF_X3 FE_OFC299_g4457A (.Z(FE_OFN299_g4457A),.A(g4457A));
BUF_X3 FE_OFC298_g3015A (.Z(FE_OFN298_g3015A),.A(FE_OFN119_g3015A));
BUF_X3 FE_OFC297_g3015A (.Z(FE_OFN297_g3015A),.A(FE_OFN348_g3015A));
INV_X1 FE_OFC296_g3914A (.ZN(FE_OFN296_g3914A),.A(FE_OFN294_g3914A));
INV_X1 FE_OFC294_g3914A (.ZN(FE_OFN294_g3914A),.A(FE_OFN113_g3914A));
BUF_X3 FE_OFC293_g3015A (.Z(FE_OFN293_g3015A),.A(FE_OFN292_g3015A));
BUF_X3 FE_OFC292_g3015A (.Z(FE_OFN292_g3015A),.A(FE_OFN345_g3015A));
BUF_X3 FE_OFC291_g4880A (.Z(FE_OFN291_g4880A),.A(FE_OFN290_g4880A));
BUF_X3 FE_OFC290_g4880A (.Z(FE_OFN290_g4880A),.A(g4880A));
BUF_X3 FE_OFC289_g4679A (.Z(FE_OFN289_g4679A),.A(g4679A));
BUF_X3 FE_OFC288_g4263A (.Z(FE_OFN288_g4263A),.A(g4263A));
INV_X1 FE_OFC287_g3586A (.ZN(FE_OFN287_g3586A),.A(FE_OFN284_g3586A));
INV_X1 FE_OFC284_g3586A (.ZN(FE_OFN284_g3586A),.A(FE_OFN110_g3586A));
BUF_X3 FE_OFC283_I8869A (.Z(FE_OFN283_I8869A),.A(FE_OFN97_I8869A));
BUF_X3 FE_OFC282_g6165A (.Z(FE_OFN282_g6165A),.A(g6165A));
BUF_X3 FE_OFC281_g2216A (.Z(FE_OFN281_g2216A),.A(FE_OFN95_g2216A));
BUF_X3 FE_OFC280_g9536A (.Z(FE_OFN280_g9536A),.A(FE_OFN64_g9536A));
BUF_X3 FE_OFC279_g11157A (.Z(FE_OFN279_g11157A),.A(g11157A));
BUF_X3 FE_OFC278_g10927A (.Z(FE_OFN278_g10927A),.A(g10927A));
BUF_X3 FE_OFC277_g48A (.Z(FE_OFN277_g48A),.A(FE_OFN276_g48A));
BUF_X3 FE_OFC276_g48A (.Z(FE_OFN276_g48A),.A(FE_OFN275_g48A));
BUF_X3 FE_OFC275_g48A (.Z(FE_OFN275_g48A),.A(g48A));
BUF_X3 FE_OFC273_g85A (.Z(FE_OFN273_g85A),.A(FE_OFN271_g85A));
BUF_X3 FE_OFC271_g85A (.Z(FE_OFN271_g85A),.A(g85A));
BUF_X3 FE_OFC269_g109A (.Z(FE_OFN269_g109A),.A(FE_OFN267_g109A));
BUF_X3 FE_OFC267_g109A (.Z(FE_OFN267_g109A),.A(g109A));
BUF_X3 FE_OFC266_g18A (.Z(FE_OFN266_g18A),.A(FE_OFN325_g18A));
BUF_X3 FE_OFC260_g18A (.Z(FE_OFN260_g18A),.A(g2355A));
BUF_X3 FE_OFC254_g461A (.Z(FE_OFN254_g461A),.A(g461A));
BUF_X3 FE_OFC253_g1786A (.Z(FE_OFN253_g1786A),.A(g1786A));
BUF_X3 FE_OFC252_g1791A (.Z(FE_OFN252_g1791A),.A(g1791A));
BUF_X3 FE_OFC251_g1801A (.Z(FE_OFN251_g1801A),.A(g1801A));
BUF_X3 FE_OFC250_g471A (.Z(FE_OFN250_g471A),.A(g471A));
BUF_X3 FE_OFC248_g466A (.Z(FE_OFN248_g466A),.A(g466A));
BUF_X3 FE_OFC247_g1771A (.Z(FE_OFN247_g1771A),.A(g1771A));
INV_X1 FE_OFC245_g1690A (.ZN(FE_OFN245_g1690A),.A(g2424A));
BUF_X3 FE_OFC241_g1690A (.Z(FE_OFN241_g1690A),.A(g1690A));
BUF_X3 FE_OFC240_g1110A (.Z(FE_OFN240_g1110A),.A(g1110A));
BUF_X3 FE_OFC239_g1796A (.Z(FE_OFN239_g1796A),.A(g1796A));
BUF_X3 FE_OFC238_g1781A (.Z(FE_OFN238_g1781A),.A(g1781A));
BUF_X3 FE_OFC237_g1806A (.Z(FE_OFN237_g1806A),.A(g1806A));
BUF_X3 FE_OFC236_g1776A (.Z(FE_OFN236_g1776A),.A(g1776A));
BUF_X3 FE_OFC235_g2024A (.Z(FE_OFN235_g2024A),.A(FE_OFN234_g2024A));
BUF_X3 FE_OFC234_g2024A (.Z(FE_OFN234_g2024A),.A(g2024A));
INV_X1 FE_OFC233_I5565A (.ZN(FE_OFN233_I5565A),.A(FE_OFN230_I5565A));
INV_X1 FE_OFC230_I5565A (.ZN(FE_OFN230_I5565A),.A(I6360A));
INV_X1 FE_OFC229_g3880A (.ZN(FE_OFN229_g3880A),.A(FE_OFN227_g3880A));
INV_X1 FE_OFC227_g3880A (.ZN(FE_OFN227_g3880A),.A(FE_OFN226_g3880A));
BUF_X3 FE_OFC226_g3880A (.Z(FE_OFN226_g3880A),.A(g3880A));
BUF_X3 FE_OFC225_g2276A (.Z(FE_OFN225_g2276A),.A(FE_OFN224_g2276A));
BUF_X3 FE_OFC224_g2276A (.Z(FE_OFN224_g2276A),.A(g2276A));
BUF_X3 FE_OFC223_g4401A (.Z(FE_OFN223_g4401A),.A(g4401A));
BUF_X3 FE_OFC221_g3440A (.Z(FE_OFN221_g3440A),.A(g3440A));
BUF_X3 FE_OFC219_g5557A (.Z(FE_OFN219_g5557A),.A(FE_OFN218_g5557A));
BUF_X3 FE_OFC218_g5557A (.Z(FE_OFN218_g5557A),.A(g5557A));
INV_X1 FE_OFC217_g5013A (.ZN(FE_OFN217_g5013A),.A(g6403A));
BUF_X3 FE_OFC213_g6003A (.Z(FE_OFN213_g6003A),.A(g6003A));
BUF_X3 FE_OFC211_g7246A (.Z(FE_OFN211_g7246A),.A(FE_OFN210_g7246A));
BUF_X3 FE_OFC210_g7246A (.Z(FE_OFN210_g7246A),.A(g7246A));
INV_X1 FE_OFC209_g6863A (.ZN(FE_OFN209_g6863A),.A(FE_OFN207_g6863A));
INV_X1 FE_OFC207_g6863A (.ZN(FE_OFN207_g6863A),.A(FE_OFN206_g6863A));
BUF_X3 FE_OFC206_g6863A (.Z(FE_OFN206_g6863A),.A(g6863A));
BUF_X3 FE_OFC204_g3664A (.Z(FE_OFN204_g3664A),.A(g3664A));
BUF_X3 FE_OFC200_g4921A (.Z(FE_OFN200_g4921A),.A(g4921A));
BUF_X3 FE_OFC199_g7697A (.Z(FE_OFN199_g7697A),.A(FE_OFN198_g7697A));
INV_X1 FE_OFC198_g7697A (.ZN(FE_OFN198_g7697A),.A(FE_OFN196_g7697A));
INV_X1 FE_OFC196_g7697A (.ZN(FE_OFN196_g7697A),.A(g7697A));
INV_X1 FE_OFC195_g6488A (.ZN(FE_OFN195_g6488A),.A(FE_OFN192_g6488A));
INV_X1 FE_OFC192_g6488A (.ZN(FE_OFN192_g6488A),.A(g6488A));
BUF_X3 FE_OFC191_g6488A (.Z(FE_OFN191_g6488A),.A(g6488A));
INV_X1 FE_OFC189_g7638A (.ZN(FE_OFN189_g7638A),.A(FE_OFN187_g7638A));
INV_X1 FE_OFC187_g7638A (.ZN(FE_OFN187_g7638A),.A(g7638A));
BUF_X3 FE_OFC184_I7048A (.Z(FE_OFN184_I7048A),.A(I7048A));
BUF_X3 FE_OFC180_g5354A (.Z(FE_OFN180_g5354A),.A(FE_OFN179_g5354A));
BUF_X3 FE_OFC179_g5354A (.Z(FE_OFN179_g5354A),.A(FE_OFN178_g5354A));
BUF_X3 FE_OFC178_g5354A (.Z(FE_OFN178_g5354A),.A(g5354A));
BUF_X3 FE_OFC177_g5919A (.Z(FE_OFN177_g5919A),.A(g5919A));
BUF_X3 FE_OFC176_g5151A (.Z(FE_OFN176_g5151A),.A(FE_OFN306_g5128A));
INV_X1 FE_OFC168_g5361A (.ZN(FE_OFN168_g5361A),.A(FE_OFN166_g5361A));
INV_X1 FE_OFC166_g5361A (.ZN(FE_OFN166_g5361A),.A(FE_OFN164_g5361A));
INV_X1 FE_OFC164_g5361A (.ZN(FE_OFN164_g5361A),.A(FE_OFN161_g5361A));
INV_X1 FE_OFC161_g5361A (.ZN(FE_OFN161_g5361A),.A(g5361A));
BUF_X3 FE_OFC160_I6424A (.Z(FE_OFN160_I6424A),.A(FE_OFN350_g3121A));
BUF_X3 FE_OFC155_g3121A (.Z(FE_OFN155_g3121A),.A(g3121A));
BUF_X3 FE_OFC154_g4640A (.Z(FE_OFN154_g4640A),.A(FE_OFN153_g4640A));
INV_X1 FE_OFC153_g4640A (.ZN(FE_OFN153_g4640A),.A(FE_OFN321_g5261A));
BUF_X4 FE_OFC147_g4682A (.Z(FE_OFN147_g4682A),.A(FE_OFN146_g4682A));
BUF_X3 FE_OFC146_g4682A (.Z(FE_OFN146_g4682A),.A(FE_OFN144_g4682A));
INV_X1 FE_OFC144_g4682A (.ZN(FE_OFN144_g4682A),.A(FE_OFN142_g4682A));
INV_X1 FE_OFC142_g4682A (.ZN(FE_OFN142_g4682A),.A(g4682A));
INV_X1 FE_OFC141_g3829A (.ZN(FE_OFN141_g3829A),.A(FE_OFN299_g4457A));
BUF_X3 FE_OFC137_g3829A (.Z(FE_OFN137_g3829A),.A(g3829A));
INV_X1 FE_OFC136_g3863A (.ZN(FE_OFN136_g3863A),.A(FE_OFN134_g3863A));
INV_X1 FE_OFC134_g3863A (.ZN(FE_OFN134_g3863A),.A(g3863A));
BUF_X3 FE_OFC133_g3015A (.Z(FE_OFN133_g3015A),.A(FE_OFN131_g3015A));
BUF_X3 FE_OFC132_g3015A (.Z(FE_OFN132_g3015A),.A(FE_OFN293_g3015A));
INV_X1 FE_OFC131_g3015A (.ZN(FE_OFN131_g3015A),.A(FE_OFN291_g4880A));
BUF_X3 FE_OFC119_g3015A (.Z(FE_OFN119_g3015A),.A(g3015A));
BUF_X3 FE_OFC118_g4807A (.Z(FE_OFN118_g4807A),.A(FE_OFN117_g4807A));
BUF_X3 FE_OFC117_g4807A (.Z(FE_OFN117_g4807A),.A(FE_OFN116_g4807A));
BUF_X3 FE_OFC116_g4807A (.Z(FE_OFN116_g4807A),.A(FE_OFN115_g4807A));
BUF_X3 FE_OFC115_g4807A (.Z(FE_OFN115_g4807A),.A(g4807A));
INV_X1 FE_OFC113_g3914A (.ZN(FE_OFN113_g3914A),.A(FE_OFN111_g3914A));
INV_X1 FE_OFC111_g3914A (.ZN(FE_OFN111_g3914A),.A(g4673A));
INV_X1 FE_OFC110_g3586A (.ZN(FE_OFN110_g3586A),.A(g4263A));
BUF_X3 FE_OFC103_g3586A (.Z(FE_OFN103_g3586A),.A(FE_OFN102_g3586A));
BUF_X3 FE_OFC102_g3586A (.Z(FE_OFN102_g3586A),.A(g3586A));
BUF_X3 FE_OFC100_g4421A (.Z(FE_OFN100_g4421A),.A(FE_OFN99_g4421A));
BUF_X3 FE_OFC99_g4421A (.Z(FE_OFN99_g4421A),.A(g4421A));
BUF_X3 FE_OFC97_I8869A (.Z(FE_OFN97_I8869A),.A(I8869A));
BUF_X3 FE_OFC96_g2169A (.Z(FE_OFN96_g2169A),.A(g2169A));
BUF_X3 FE_OFC95_g2216A (.Z(FE_OFN95_g2216A),.A(FE_OFN93_g2216A));
BUF_X3 FE_OFC93_g2216A (.Z(FE_OFN93_g2216A),.A(FE_OFN92_g2216A));
BUF_X3 FE_OFC92_g2216A (.Z(FE_OFN92_g2216A),.A(g2216A));
BUF_X3 FE_OFC91_g2172A (.Z(FE_OFN91_g2172A),.A(g2172A));
BUF_X3 FE_OFC90_I11360A (.Z(FE_OFN90_I11360A),.A(FE_OFN89_I11360A));
BUF_X3 FE_OFC89_I11360A (.Z(FE_OFN89_I11360A),.A(I11360A));
BUF_X3 FE_OFC88_g2178A (.Z(FE_OFN88_g2178A),.A(g2178A));
BUF_X3 FE_OFC87_g2176A (.Z(FE_OFN87_g2176A),.A(FE_OFN86_g2176A));
BUF_X3 FE_OFC86_g2176A (.Z(FE_OFN86_g2176A),.A(FE_OFN85_g2176A));
BUF_X3 FE_OFC85_g2176A (.Z(FE_OFN85_g2176A),.A(FE_OFN83_g2176A));
INV_X1 FE_OFC84_g2176A (.ZN(FE_OFN84_g2176A),.A(FE_OFN81_g2176A));
INV_X1 FE_OFC83_g2176A (.ZN(FE_OFN83_g2176A),.A(FE_OFN81_g2176A));
INV_X1 FE_OFC82_g2176A (.ZN(FE_OFN82_g2176A),.A(FE_OFN81_g2176A));
INV_X1 FE_OFC81_g2176A (.ZN(FE_OFN81_g2176A),.A(g2176A));
BUF_X3 FE_OFC80_g2175A (.Z(FE_OFN80_g2175A),.A(g2175A));
INV_X1 FE_OFC79_g8700A (.ZN(FE_OFN79_g8700A),.A(g9097A));
BUF_X3 FE_OFC76_g8700A (.Z(FE_OFN76_g8700A),.A(g8700A));
BUF_X3 FE_OFC73_g8858A (.Z(FE_OFN73_g8858A),.A(g8858A));
BUF_X3 FE_OFC72_g9292A (.Z(FE_OFN72_g9292A),.A(FE_OFN71_g9292A));
BUF_X3 FE_OFC71_g9292A (.Z(FE_OFN71_g9292A),.A(g9292A));
BUF_X3 FE_OFC70_g9490A (.Z(FE_OFN70_g9490A),.A(g9490A));
BUF_X3 FE_OFC69_g9392A (.Z(FE_OFN69_g9392A),.A(FE_OFN68_g9392A));
BUF_X3 FE_OFC68_g9392A (.Z(FE_OFN68_g9392A),.A(g9392A));
BUF_X3 FE_OFC67_g9367A (.Z(FE_OFN67_g9367A),.A(g9367A));
BUF_X3 FE_OFC64_g9536A (.Z(FE_OFN64_g9536A),.A(g9536A));
BUF_X3 FE_OFC63_g9474A (.Z(FE_OFN63_g9474A),.A(g9474A));
BUF_X3 FE_OFC62_g9274A (.Z(FE_OFN62_g9274A),.A(g9274A));
BUF_X3 FE_OFC61_g9624A (.Z(FE_OFN61_g9624A),.A(FE_OFN60_g9624A));
BUF_X3 FE_OFC60_g9624A (.Z(FE_OFN60_g9624A),.A(g9624A));
INV_X1 FE_OFC59_g9432A (.ZN(FE_OFN59_g9432A),.A(FE_OFN57_g9432A));
INV_X1 FE_OFC57_g9432A (.ZN(FE_OFN57_g9432A),.A(g9432A));
BUF_X3 FE_OFC56_g9052A (.Z(FE_OFN56_g9052A),.A(FE_OFN54_g9052A));
BUF_X3 FE_OFC54_g9052A (.Z(FE_OFN54_g9052A),.A(g9052A));
BUF_X3 FE_OFC53_g9173A (.Z(FE_OFN53_g9173A),.A(FE_OFN52_g9173A));
BUF_X3 FE_OFC52_g9173A (.Z(FE_OFN52_g9173A),.A(g9173A));
BUF_X3 FE_OFC51_g9111A (.Z(FE_OFN51_g9111A),.A(g9111A));
BUF_X3 FE_OFC50_g9030A (.Z(FE_OFN50_g9030A),.A(FE_OFN49_g9030A));
BUF_X3 FE_OFC49_g9030A (.Z(FE_OFN49_g9030A),.A(g9030A));
BUF_X3 FE_OFC48_g9151A (.Z(FE_OFN48_g9151A),.A(FE_OFN47_g9151A));
BUF_X3 FE_OFC47_g9151A (.Z(FE_OFN47_g9151A),.A(g9151A));
BUF_X3 FE_OFC46_g9125A (.Z(FE_OFN46_g9125A),.A(FE_OFN45_g9125A));
BUF_X3 FE_OFC45_g9125A (.Z(FE_OFN45_g9125A),.A(FE_OFN44_g9125A));
BUF_X3 FE_OFC44_g9125A (.Z(FE_OFN44_g9125A),.A(g9125A));
BUF_X3 FE_OFC42_g9205A (.Z(FE_OFN42_g9205A),.A(g9205A));
BUF_X3 FE_OFC40_g9240A (.Z(FE_OFN40_g9240A),.A(g9240A));
BUF_X3 FE_OFC39_g9223A (.Z(FE_OFN39_g9223A),.A(g9223A));
BUF_X3 FE_OFC35_g9785A (.Z(FE_OFN35_g9785A),.A(FE_OFN34_g9785A));
BUF_X3 FE_OFC34_g9785A (.Z(FE_OFN34_g9785A),.A(g9785A));
BUF_X3 FE_OFC33_g9454A (.Z(FE_OFN33_g9454A),.A(FE_OFN32_g9454A));
BUF_X3 FE_OFC32_g9454A (.Z(FE_OFN32_g9454A),.A(g9454A));
BUF_X3 FE_OFC27_g11519A (.Z(FE_OFN27_g11519A),.A(g11519A));
BUF_X3 FE_OFC21_g10702A (.Z(FE_OFN21_g10702A),.A(FE_OFN20_g10702A));
BUF_X3 FE_OFC20_g10702A (.Z(FE_OFN20_g10702A),.A(FE_OFN18_g10702A));
BUF_X3 FE_OFC18_g10702A (.Z(FE_OFN18_g10702A),.A(FE_OFN13_g10702A));
INV_X1 FE_OFC17_g10702A (.ZN(FE_OFN17_g10702A),.A(FE_OFN15_g10702A));
INV_X1 FE_OFC15_g10702A (.ZN(FE_OFN15_g10702A),.A(FE_OFN14_g10702A));
BUF_X3 FE_OFC14_g10702A (.Z(FE_OFN14_g10702A),.A(FE_OFN9_g10702A));
INV_X1 FE_OFC13_g10702A (.ZN(FE_OFN13_g10702A),.A(FE_OFN10_g10702A));
INV_X1 FE_OFC10_g10702A (.ZN(FE_OFN10_g10702A),.A(FE_OFN9_g10702A));
BUF_X3 FE_OFC9_g10702A (.Z(FE_OFN9_g10702A),.A(FE_OFN8_g10702A));
BUF_X3 FE_OFC8_g10702A (.Z(FE_OFN8_g10702A),.A(FE_OFN7_g10702A));
BUF_X3 FE_OFC7_g10702A (.Z(FE_OFN7_g10702A),.A(g10702A));
BUF_X3 FE_OFC4_g10950A (.Z(FE_OFN4_g10950A),.A(FE_OFN3_g10950A));
INV_X1 FE_OFC3_g10950A (.ZN(FE_OFN3_g10950A),.A(FE_OFN0_g10950A));
INV_X1 FE_OFC0_g10950A (.ZN(FE_OFN0_g10950A),.A(g10950A));
INV_X1 U_g2299A (.ZN(g2299A),.A(g1707A));
INV_X1 U_g9291A (.ZN(g9291A),.A(FE_OFN79_g8700A));
INV_X4 U_I7048A (.ZN(I7048A),.A(g2807A));
INV_X1 U_g1981A (.ZN(g1981A),.A(g650A));
INV_X1 U_g3982A (.ZN(g3982A),.A(g2118A));
INV_X1 U_g3629A (.ZN(g3629A),.A(FE_OFN266_g18A));
INV_X1 U_g6842A (.ZN(g6842A),.A(I9769A));
INV_X1 U_g8617A (.ZN(g8617A),.A(g8465A));
INV_X1 U_g2078A (.ZN(g2078A),.A(g135A));
INV_X1 U_g2340A (.ZN(g2340A),.A(g1918A));
INV_X1 U_g7684A (.ZN(g7684A),.A(FE_OFN83_g2176A));
INV_X1 U_g3800A (.ZN(g3800A),.A(FE_OFN250_g471A));
INV_X1 U_g6941A (.ZN(g6941A),.A(FE_OFN88_g2178A));
INV_X1 U_g2435A (.ZN(g2435A),.A(g201A));
INV_X4 U_g4010A (.ZN(g4010A),.A(g3744A));
INV_X1 U_g2082A (.ZN(g2082A),.A(g1371A));
INV_X1 U_g5519A (.ZN(g5519A),.A(g4811A));
INV_X1 U_g10668A (.ZN(g10668A),.A(g10563A));
INV_X1 U_g4172A (.ZN(g4172A),.A(g2057A));
INV_X1 U_g8709A (.ZN(g8709A),.A(g8451A));
INV_X1 U_g2214A (.ZN(g2214A),.A(g115A));
INV_X1 U_I7847A (.ZN(I7847A),.A(g3435A));
INV_X1 U_g8340A (.ZN(g8340A),.A(I13400A));
INV_X1 U_g4566A (.ZN(g4566A),.A(g3753A));
INV_X1 U_g3348A (.ZN(g3348A),.A(FE_OFN267_g109A));
INV_X1 U_I15968A (.ZN(I15968A),.A(g10408A));
INV_X1 U_g11060A (.ZN(g11060A),.A(g10937A));
INV_X1 U_I15855A (.ZN(I15855A),.A(g10336A));
INV_X1 U_g6270A (.ZN(g6270A),.A(I9383A));
INV_X1 U_g10679A (.ZN(g10679A),.A(g10584A));
INV_X1 U_g1968A (.ZN(g1968A),.A(g369A));
INV_X1 U_g5659A (.ZN(g5659A),.A(I7771A));
INV_X1 U_I15503A (.ZN(I15503A),.A(g9995A));
INV_X1 U_g8110A (.ZN(g8110A),.A(g7996A));
INV_X1 U_g2556A (.ZN(g2556A),.A(g186A));
INV_X1 U_I7817A (.ZN(I7817A),.A(g3399A));
INV_X1 U_g2222A (.ZN(g2222A),.A(g158A));
INV_X1 U_I13373A (.ZN(I13373A),.A(g8226A));
INV_X1 U_g4202A (.ZN(g4202A),.A(I5430A));
INV_X1 U_I9880A (.ZN(I9880A),.A(g5405A));
INV_X1 U_g4094A (.ZN(g4094A),.A(g2744A));
INV_X1 U_g4567A (.ZN(g4567A),.A(g3374A));
INV_X1 U_I14312A (.ZN(I14312A),.A(g8814A));
INV_X1 U_g11111A (.ZN(g11111A),.A(g10702A));
INV_X1 U_g4776A (.ZN(g4776A),.A(FE_OFN344_g3586A));
INV_X1 U_I15986A (.ZN(I15986A),.A(g10417A));
INV_X1 U_g2237A (.ZN(g2237A),.A(g713A));
INV_X1 U_g7897A (.ZN(g7897A),.A(g7712A));
INV_X1 U_g3121A (.ZN(g3121A),.A(FE_OFN352_g109A));
INV_X1 U_g5420A (.ZN(g5420A),.A(g4300A));
INV_X1 U_g10455A (.ZN(g10455A),.A(I15956A));
INV_X1 U_g2557A (.ZN(g2557A),.A(g1840A));
INV_X1 U_g9097A (.ZN(g9097A),.A(g8700A));
INV_X1 U_g3938A (.ZN(g3938A),.A(g2299A));
INV_X1 U_g8563A (.ZN(g8563A),.A(I7829A));
INV_X1 U_g6259A (.ZN(g6259A),.A(g2175A));
INV_X1 U_g4179A (.ZN(g4179A),.A(g1992A));
INV_X1 U_g7682A (.ZN(g7682A),.A(FE_OFN83_g2176A));
INV_X1 U_g4379A (.ZN(g4379A),.A(g3698A));
INV_X1 U_I4917A (.ZN(I4917A),.A(g584A));
INV_X1 U_g2254A (.ZN(g2254A),.A(g131A));
INV_X1 U_g4289A (.ZN(g4289A),.A(FE_OFN298_g3015A));
INV_X1 U_g4777A (.ZN(g4777A),.A(g3992A));
INV_X1 U_g8089A (.ZN(g8089A),.A(g7934A));
INV_X1 U_g2438A (.ZN(g2438A),.A(g243A));
INV_X1 U_g4271A (.ZN(g4271A),.A(g2024A));
INV_X1 U_g7045A (.ZN(g7045A),.A(g6003A));
INV_X1 U_I5424A (.ZN(I5424A),.A(g910A));
INV_X1 U_g2212A (.ZN(g2212A),.A(g686A));
INV_X1 U_g3141A (.ZN(g3141A),.A(g2563A));
INV_X1 U_g3710A (.ZN(g3710A),.A(g3215A));
INV_X1 U_g7920A (.ZN(g7920A),.A(g7516A));
INV_X1 U_g2229A (.ZN(g2229A),.A(g162A));
INV_X1 U_I15157A (.ZN(I15157A),.A(g9931A));
INV_X1 U_g11157A (.ZN(g11157A),.A(FE_OFN3_g10950A));
INV_X1 U_g4209A (.ZN(g4209A),.A(I5002A));
INV_X1 U_I9279A (.ZN(I9279A),.A(g91A));
INV_X1 U_I5044A (.ZN(I5044A),.A(g1182A));
INV_X1 U_I15287A (.ZN(I15287A),.A(g9968A));
INV_X1 U_g2249A (.ZN(g2249A),.A(g127A));
INV_X1 U_g11596A (.ZN(g11596A),.A(g11580A));
INV_X1 U_g11243A (.ZN(g11243A),.A(FE_OFN8_g10702A));
INV_X1 U_g6266A (.ZN(g6266A),.A(g2208A));
INV_X1 U_g8062A (.ZN(g8062A),.A(I4783A));
INV_X1 U_I5414A (.ZN(I5414A),.A(g904A));
INV_X1 U_g3628A (.ZN(g3628A),.A(g3111A));
INV_X1 U_g6255A (.ZN(g6255A),.A(I9237A));
INV_X1 U_g4175A (.ZN(g4175A),.A(g1988A));
INV_X1 U_g6081A (.ZN(g6081A),.A(g4977A));
INV_X1 U_g7910A (.ZN(g7910A),.A(g7460A));
INV_X1 U_g4285A (.ZN(g4285A),.A(g3688A));
INV_X1 U_g6354A (.ZN(g6354A),.A(g5867A));
INV_X1 U_g2031A (.ZN(g2031A),.A(g1690A));
INV_X1 U_g8085A (.ZN(g8085A),.A(g7932A));
INV_X1 U_g2176A (.ZN(g2176A),.A(g82A));
INV_X1 U_g7883A (.ZN(g7883A),.A(g7246A));
INV_X1 U_g4737A (.ZN(g4737A),.A(g3440A));
INV_X1 U_I13351A (.ZN(I13351A),.A(g8214A));
INV_X1 U_g6267A (.ZN(g6267A),.A(I9326A));
INV_X1 U_g3440A (.ZN(g3440A),.A(g3041A));
INV_X1 U_g2610A (.ZN(g2610A),.A(I4917A));
INV_X1 U_g4205A (.ZN(g4205A),.A(I4992A));
INV_X1 U_g10883A (.ZN(g10883A),.A(g10809A));
INV_X1 U_g5521A (.ZN(g5521A),.A(FE_OFN221_g3440A));
INV_X1 U_I6260A (.ZN(I6260A),.A(g1696A));
INV_X1 U_I9311A (.ZN(I9311A),.A(g103A));
INV_X1 U_I5579A (.ZN(I5579A),.A(g1197A));
INV_X1 U_g10439A (.ZN(g10439A),.A(g10334A));
INV_X1 U_g5878A (.ZN(g5878A),.A(g5309A));
INV_X1 U_g6932A (.ZN(g6932A),.A(I7829A));
INV_X1 U_g4273A (.ZN(g4273A),.A(FE_OFN133_g3015A));
INV_X1 U_g5658A (.ZN(g5658A),.A(I7752A));
INV_X1 U_g7467A (.ZN(g7467A),.A(FE_OFN84_g2176A));
INV_X1 U_g1990A (.ZN(g1990A),.A(g774A));
INV_X1 U_I13436A (.ZN(I13436A),.A(g8187A));
INV_X1 U_g2399A (.ZN(g2399A),.A(g605A));
INV_X1 U_g8980A (.ZN(g8980A),.A(I14306A));
INV_X1 U_g6716A (.ZN(g6716A),.A(FE_OFN115_g4807A));
INV_X1 U_g7685A (.ZN(g7685A),.A(FE_OFN87_g2176A));
INV_X1 U_g8849A (.ZN(g8849A),.A(g8745A));
INV_X1 U_I7840A (.ZN(I7840A),.A(g3431A));
INV_X1 U_g10852A (.ZN(g10852A),.A(g10739A));
INV_X1 U_g7562A (.ZN(g7562A),.A(FE_OFN91_g2172A));
INV_X1 U_g6258A (.ZN(g6258A),.A(g2172A));
INV_X1 U_g4178A (.ZN(g4178A),.A(g1991A));
INV_X4 U_g4679A (.ZN(g4679A),.A(FE_OFN293_g3015A));
INV_X1 U_g3776A (.ZN(g3776A),.A(g2579A));
INV_X1 U_g2008A (.ZN(g2008A),.A(g971A));
INV_X1 U_g6274A (.ZN(g6274A),.A(I9293A));
INV_X1 U_g2336A (.ZN(g2336A),.A(g1900A));
INV_X1 U_g3521A (.ZN(g3521A),.A(FE_OFN359_g18A));
INV_X1 U_g6280A (.ZN(g6280A),.A(g2253A));
INV_X1 U_I6962A (.ZN(I6962A),.A(g2791A));
INV_X1 U_g2230A (.ZN(g2230A),.A(g704A));
INV_X1 U_g4437A (.ZN(g4437A),.A(FE_OFN235_g2024A));
INV_X1 U_g4208A (.ZN(g4208A),.A(I5588A));
INV_X1 U_g7505A (.ZN(g7505A),.A(FE_OFN87_g2176A));
INV_X1 U_I15974A (.ZN(I15974A),.A(g10411A));
INV_X1 U_g2550A (.ZN(g2550A),.A(g1834A));
INV_X1 U_g10400A (.ZN(g10400A),.A(g10348A));
INV_X1 U_I9282A (.ZN(I9282A),.A(g101A));
INV_X1 U_I5584A (.ZN(I5584A),.A(g1200A));
INV_X4 U_g9490A (.ZN(g9490A),.A(g9324A));
INV_X1 U_g2395A (.ZN(g2395A),.A(g231A));
INV_X1 U_g8465A (.ZN(g8465A),.A(g8289A));
INV_X1 U_g6403A (.ZN(g6403A),.A(g5013A));
INV_X1 U_I15510A (.ZN(I15510A),.A(g10013A));
INV_X1 U_g2248A (.ZN(g2248A),.A(g99A));
INV_X1 U_g3744A (.ZN(g3744A),.A(FE_OFN269_g109A));
INV_X1 U_I4883A (.ZN(I4883A),.A(g581A));
INV_X1 U_g7688A (.ZN(g7688A),.A(FE_OFN83_g2176A));
INV_X1 U_g2481A (.ZN(g2481A),.A(g882A));
INV_X1 U_g10683A (.ZN(g10683A),.A(g10385A));
INV_X1 U_I5070A (.ZN(I5070A),.A(g1194A));
INV_X1 U_g4888A (.ZN(g4888A),.A(I5101A));
INV_X1 U_g4171A (.ZN(g4171A),.A(I6962A));
INV_X1 U_g4787A (.ZN(g4787A),.A(g3423A));
INV_X1 U_g6447A (.ZN(g6447A),.A(FE_OFN218_g5557A));
INV_X1 U_g3092A (.ZN(g3092A),.A(g639A));
INV_X1 U_g4281A (.ZN(g4281A),.A(g3586A));
INV_X1 U_g5613A (.ZN(g5613A),.A(FE_OFN131_g3015A));
INV_X1 U_g8255A (.ZN(g8255A),.A(g7986A));
INV_X1 U_g8081A (.ZN(g8081A),.A(g8000A));
INV_X1 U_I5406A (.ZN(I5406A),.A(g898A));
INV_X1 U_I4780A (.ZN(I4780A),.A(g872A));
INV_X1 U_g10584A (.ZN(g10584A),.A(g10522A));
INV_X1 U_g6272A (.ZN(g6272A),.A(I9268A));
INV_X1 U_g8783A (.ZN(g8783A),.A(g8746A));
INV_X1 U_g8979A (.ZN(g8979A),.A(I14303A));
INV_X1 U_g4201A (.ZN(g4201A),.A(I5427A));
INV_X1 U_I5445A (.ZN(I5445A),.A(g922A));
INV_X1 U_g4449A (.ZN(g4449A),.A(g4144A));
INV_X1 U_g7696A (.ZN(g7696A),.A(FE_OFN86_g2176A));
INV_X1 U_g8828A (.ZN(g8828A),.A(g8744A));
INV_X1 U_g2677A (.ZN(g2677A),.A(g2034A));
INV_X1 U_g10361A (.ZN(g10361A),.A(g10268A));
INV_X1 U_g3737A (.ZN(g3737A),.A(g2506A));
INV_X1 U_I9332A (.ZN(I9332A),.A(g104A));
INV_X1 U_g9525A (.ZN(g9525A),.A(g9257A));
INV_X1 U_g2198A (.ZN(g2198A),.A(g668A));
INV_X1 U_I7771A (.ZN(I7771A),.A(g3418A));
INV_X1 U_g3523A (.ZN(g3523A),.A(g1845A));
INV_X1 U_g2241A (.ZN(g2241A),.A(g722A));
INV_X1 U_g7681A (.ZN(g7681A),.A(FE_OFN87_g2176A));
INV_X1 U_g7697A (.ZN(g7697A),.A(g7101A));
INV_X1 U_g7914A (.ZN(g7914A),.A(g7651A));
INV_X1 U_g8349A (.ZN(g8349A),.A(I13427A));
INV_X1 U_g6260A (.ZN(g6260A),.A(g2178A));
INV_X1 U_I14319A (.ZN(I14319A),.A(g8816A));
INV_X1 U_g10463A (.ZN(g10463A),.A(I15980A));
INV_X1 U_I5388A (.ZN(I5388A),.A(g889A));
INV_X1 U_g2211A (.ZN(g2211A),.A(g153A));
INV_X1 U_g6279A (.ZN(g6279A),.A(g2248A));
INV_X1 U_g3983A (.ZN(g3983A),.A(g3222A));
INV_X1 U_I5430A (.ZN(I5430A),.A(g916A));
INV_X4 U_g4678A (.ZN(g4678A),.A(g3546A));
INV_X1 U_g3543A (.ZN(g3543A),.A(g3101A));
INV_X1 U_g9507A (.ZN(g9507A),.A(g9268A));
INV_X1 U_g10421A (.ZN(g10421A),.A(g10331A));
INV_X1 U_g8352A (.ZN(g8352A),.A(I13436A));
INV_X1 U_g7460A (.ZN(g7460A),.A(FE_OFN85_g2176A));
INV_X1 U_g2083A (.ZN(g2083A),.A(g139A));
INV_X1 U_I6360A (.ZN(I6360A),.A(g1713A));
INV_X1 U_I4992A (.ZN(I4992A),.A(g1170A));
INV_X1 U_I16982A (.ZN(I16982A),.A(g10629A));
INV_X1 U_g8599A (.ZN(g8599A),.A(g8546A));
INV_X1 U_g6253A (.ZN(g6253A),.A(I9479A));
INV_X1 U_g2061A (.ZN(g2061A),.A(g1828A));
INV_X1 U_g2187A (.ZN(g2187A),.A(g746A));
INV_X1 U_g4173A (.ZN(g4173A),.A(g1984A));
INV_X1 U_g8984A (.ZN(g8984A),.A(I14319A));
INV_X1 U_g2446A (.ZN(g2446A),.A(g1400A));
INV_X1 U_g11575A (.ZN(g11575A),.A(g11561A));
INV_X1 U_g2345A (.ZN(g2345A),.A(g1936A));
INV_X1 U_g8106A (.ZN(g8106A),.A(g7950A));
INV_X1 U_g6586A (.ZN(g6586A),.A(FE_OFN118_g4807A));
INV_X1 U_g8061A (.ZN(g8061A),.A(I4780A));
INV_X1 U_g5808A (.ZN(g5808A),.A(g85A));
INV_X1 U_I5418A (.ZN(I5418A),.A(g907A));
INV_X1 U_g4203A (.ZN(g4203A),.A(I5441A));
INV_X1 U_g2016A (.ZN(g2016A),.A(g1361A));
INV_X1 U_I16252A (.ZN(I16252A),.A(g10515A));
INV_X1 U_I9273A (.ZN(I9273A),.A(g47A));
INV_X1 U_g2251A (.ZN(g2251A),.A(g731A));
INV_X1 U_g2047A (.ZN(g2047A),.A(g1857A));
INV_X1 U_g10927A (.ZN(g10927A),.A(FE_OFN17_g10702A));
INV_X1 U_g6275A (.ZN(g6275A),.A(I9308A));
INV_X1 U_g4216A (.ZN(g4216A),.A(I5070A));
INV_X1 U_g8858A (.ZN(g8858A),.A(g8743A));
INV_X1 U_g4671A (.ZN(g4671A),.A(g3354A));
INV_X1 U_g8115A (.ZN(g8115A),.A(g7953A));
INV_X1 U_g2612A (.ZN(g2612A),.A(I4948A));
INV_X1 U_g2017A (.ZN(g2017A),.A(g1218A));
INV_X1 U_g6284A (.ZN(g6284A),.A(I9332A));
INV_X1 U_g7683A (.ZN(g7683A),.A(FE_OFN87_g2176A));
INV_X1 U_I5101A (.ZN(I5101A),.A(g1960A));
INV_X1 U_g2328A (.ZN(g2328A),.A(g1882A));
INV_X1 U_g2542A (.ZN(g2542A),.A(g1868A));
INV_X1 U_g2330A (.ZN(g2330A),.A(g1891A));
INV_X1 U_g7949A (.ZN(g7949A),.A(FE_OFN211_g7246A));
INV_X1 U_I5041A (.ZN(I5041A),.A(g1179A));
INV_X1 U_g1992A (.ZN(g1992A),.A(g782A));
INV_X1 U_g8978A (.ZN(g8978A),.A(I14299A));
INV_X1 U_I5441A (.ZN(I5441A),.A(g919A));
INV_X1 U_g4365A (.ZN(g4365A),.A(g3880A));
INV_X1 U_g8982A (.ZN(g8982A),.A(I14312A));
INV_X1 U_g8234A (.ZN(g8234A),.A(FE_OFN198_g7697A));
INV_X1 U_g8328A (.ZN(g8328A),.A(I13364A));
INV_X1 U_g4196A (.ZN(g4196A),.A(I5245A));
INV_X1 U_g2456A (.ZN(g2456A),.A(g1397A));
INV_X1 U_g7919A (.ZN(g7919A),.A(g7512A));
INV_X1 U_g5105A (.ZN(g5105A),.A(I4783A));
INV_X1 U_g1976A (.ZN(g1976A),.A(g643A));
INV_X1 U_g7952A (.ZN(g7952A),.A(FE_OFN210_g7246A));
INV_X1 U_I4820A (.ZN(I4820A),.A(g865A));
INV_X1 U_g2355A (.ZN(g2355A),.A(I5435A));
INV_X1 U_I14315A (.ZN(I14315A),.A(g8815A));
INV_X1 U_g4467A (.ZN(g4467A),.A(g3829A));
INV_X1 U_g4290A (.ZN(g4290A),.A(FE_OFN102_g3586A));
INV_X1 U_g7527A (.ZN(g7527A),.A(FE_OFN85_g2176A));
INV_X1 U_I9265A (.ZN(I9265A),.A(g46A));
INV_X1 U_g8056A (.ZN(g8056A),.A(g7671A));
INV_X1 U_g4181A (.ZN(g4181A),.A(g2449A));
INV_X1 U_g4381A (.ZN(g4381A),.A(FE_OFN296_g3914A));
INV_X1 U_g2118A (.ZN(g2118A),.A(g1854A));
INV_X1 U_I6273A (.ZN(I6273A),.A(FE_OFN363_I5565A));
INV_X1 U_g10629A (.ZN(g10629A),.A(g10583A));
INV_X1 U_g4197A (.ZN(g4197A),.A(I5410A));
INV_X1 U_g2652A (.ZN(g2652A),.A(g2008A));
INV_X1 U_g2057A (.ZN(g2057A),.A(g754A));
INV_X1 U_g10628A (.ZN(g10628A),.A(I16252A));
INV_X1 U_g3539A (.ZN(g3539A),.A(g3015A));
INV_X1 U_g4263A (.ZN(g4263A),.A(FE_OFN103_g3586A));
INV_X1 U_I9296A (.ZN(I9296A),.A(g102A));
INV_X1 U_I13323A (.ZN(I13323A),.A(g8203A));
INV_X1 U_g2549A (.ZN(g2549A),.A(g1386A));
INV_X1 U_g6278A (.ZN(g6278A),.A(I9371A));
INV_X1 U_g5261A (.ZN(g5261A),.A(g4640A));
INV_X1 U_g3419A (.ZN(g3419A),.A(g3104A));
INV_X1 U_I7829A (.ZN(I7829A),.A(g3425A));
INV_X1 U_g7516A (.ZN(g7516A),.A(FE_OFN82_g2176A));
INV_X1 U_g6282A (.ZN(g6282A),.A(I9296A));
INV_X1 U_g9802A (.ZN(g9802A),.A(g9490A));
INV_X1 U_g8318A (.ZN(g8318A),.A(I13338A));
INV_X1 U_g3086A (.ZN(g3086A),.A(g2276A));
INV_X1 U_g2253A (.ZN(g2253A),.A(g100A));
INV_X1 U_I9371A (.ZN(I9371A),.A(g96A));
INV_X1 U_I5383A (.ZN(I5383A),.A(g886A));
INV_X1 U_g2606A (.ZN(g2606A),.A(I4876A));
INV_X1 U_I5588A (.ZN(I5588A),.A(g1203A));
INV_X1 U_g7907A (.ZN(g7907A),.A(g7664A));
INV_X1 U_g4673A (.ZN(g4673A),.A(FE_OFN348_g3015A));
INV_X1 U_g2570A (.ZN(g2570A),.A(g207A));
INV_X1 U_g7915A (.ZN(g7915A),.A(g7473A));
INV_X1 U_g10377A (.ZN(g10377A),.A(I15855A));
INV_X1 U_g6264A (.ZN(g6264A),.A(g2176A));
INV_X1 U_g2607A (.ZN(g2607A),.A(I4883A));
INV_X1 U_g2506A (.ZN(g2506A),.A(g636A));
INV_X1 U_I16717A (.ZN(I16717A),.A(g10779A));
INV_X1 U_g3491A (.ZN(g3491A),.A(g1107A));
INV_X1 U_I7852A (.ZN(I7852A),.A(g3438A));
INV_X1 U_g2275A (.ZN(g2275A),.A(g757A));
INV_X1 U_g3007A (.ZN(g3007A),.A(I6240A));
INV_X1 U_g2374A (.ZN(g2374A),.A(g591A));
INV_X1 U_I9268A (.ZN(I9268A),.A(g90A));
INV_X1 U_g9424A (.ZN(g9424A),.A(g9291A));
INV_X1 U_g6271A (.ZN(g6271A),.A(I9259A));
INV_X1 U_g3793A (.ZN(g3793A),.A(FE_OFN248_g466A));
INV_X1 U_I7825A (.ZN(I7825A),.A(g3414A));
INV_X1 U_g2420A (.ZN(g2420A),.A(g237A));
INV_X1 U_g3664A (.ZN(g3664A),.A(g3209A));
INV_X1 U_g5509A (.ZN(g5509A),.A(g4739A));
INV_X1 U_g8985A (.ZN(g8985A),.A(I14326A));
INV_X1 U_g4608A (.ZN(g4608A),.A(FE_OFN141_g3829A));
INV_X1 U_g5816A (.ZN(g5816A),.A(g1810A));
INV_X1 U_I5060A (.ZN(I5060A),.A(g1191A));
INV_X1 U_I14306A (.ZN(I14306A),.A(g8812A));
INV_X1 U_g9961A (.ZN(g9961A),.A(I15157A));
INV_X1 U_g7438A (.ZN(g7438A),.A(FE_OFN195_g6488A));
INV_X1 U_g8100A (.ZN(g8100A),.A(g7947A));
INV_X1 U_g5101A (.ZN(g5101A),.A(I4780A));
INV_X1 U_g7918A (.ZN(g7918A),.A(g7505A));
INV_X1 U_g6262A (.ZN(g6262A),.A(I9273A));
INV_X1 U_g2648A (.ZN(g2648A),.A(I4820A));
INV_X1 U_g2410A (.ZN(g2410A),.A(g1453A));
INV_X1 U_g8323A (.ZN(g8323A),.A(I13351A));
INV_X1 U_I5053A (.ZN(I5053A),.A(g1188A));
INV_X1 U_g6285A (.ZN(g6285A),.A(I9352A));
INV_X1 U_g2172A (.ZN(g2172A),.A(g43A));
INV_X1 U_I13364A (.ZN(I13364A),.A(g8221A));
INV_X1 U_g2343A (.ZN(g2343A),.A(g1927A));
INV_X1 U_g4210A (.ZN(g4210A),.A(I5020A));
INV_X1 U_I4876A (.ZN(I4876A),.A(g580A));
INV_X1 U_g8566A (.ZN(g8566A),.A(I7852A));
INV_X1 U_g2202A (.ZN(g2202A),.A(g148A));
INV_X1 U_g6926A (.ZN(g6926A),.A(I7825A));
INV_X1 U_g8548A (.ZN(g8548A),.A(g8390A));
INV_X1 U_g2518A (.ZN(g2518A),.A(g590A));
INV_X1 U_g6273A (.ZN(g6273A),.A(I9279A));
INV_X1 U_g10801A (.ZN(g10801A),.A(I16507A));
INV_X1 U_g4739A (.ZN(g4739A),.A(g4117A));
INV_X1 U_g6269A (.ZN(g6269A),.A(I9368A));
INV_X1 U_g8313A (.ZN(g8313A),.A(I13323A));
INV_X1 U_I9308A (.ZN(I9308A),.A(g93A));
INV_X1 U_g4294A (.ZN(g4294A),.A(g3664A));
INV_X1 U_g3723A (.ZN(g3723A),.A(g3071A));
INV_X1 U_g10457A (.ZN(g10457A),.A(I15962A));
INV_X1 U_g8094A (.ZN(g8094A),.A(g7987A));
INV_X1 U_g2050A (.ZN(g2050A),.A(g1861A));
INV_X1 U_g7473A (.ZN(g7473A),.A(FE_OFN87_g2176A));
INV_X1 U_g2777A (.ZN(g2777A),.A(FE_OFN224_g2276A));
INV_X1 U_g2271A (.ZN(g2271A),.A(g877A));
INV_X1 U_g2611A (.ZN(g2611A),.A(I4935A));
INV_X1 U_g3368A (.ZN(g3368A),.A(g2459A));
INV_X1 U_g1987A (.ZN(g1987A),.A(g762A));
INV_X4 U_I8869A (.ZN(I8869A),.A(g4421A));
INV_X1 U_I9290A (.ZN(I9290A),.A(FE_OFN277_g48A));
INV_X1 U_I4948A (.ZN(I4948A),.A(g586A));
INV_X1 U_g8271A (.ZN(g8271A),.A(g1810A));
INV_X1 U_g1991A (.ZN(g1991A),.A(g778A));
INV_X1 U_g11199A (.ZN(g11199A),.A(FE_OFN21_g10702A));
INV_X1 U_g8981A (.ZN(g8981A),.A(I14309A));
INV_X1 U_I15365A (.ZN(I15365A),.A(g10025A));
INV_X1 U_g7852A (.ZN(g7852A),.A(FE_OFN209_g6863A));
INV_X1 U_g7923A (.ZN(g7923A),.A(g7527A));
INV_X1 U_g10431A (.ZN(g10431A),.A(g10328A));
INV_X1 U_g6265A (.ZN(g6265A),.A(I9276A));
INV_X1 U_g4782A (.ZN(g4782A),.A(g4089A));
INV_X1 U_g4292A (.ZN(g4292A),.A(FE_OFN136_g3863A));
INV_X1 U_g3760A (.ZN(g3760A),.A(g3003A));
INV_X1 U_I5435A (.ZN(I5435A),.A(g18A));
INV_X1 U_g5117A (.ZN(g5117A),.A(FE_OFN144_g4682A));
INV_X4 U_g2175A (.ZN(g2175A),.A(g44A));
INV_X1 U_I9368A (.ZN(I9368A),.A(g87A));
INV_X4 U_g2024A (.ZN(g2024A),.A(g1718A));
INV_X1 U_g6281A (.ZN(g6281A),.A(I9282A));
INV_X1 U_g3327A (.ZN(g3327A),.A(g23A));
INV_X4 U_g2424A (.ZN(g2424A),.A(FE_OFN241_g1690A));
INV_X1 U_I5002A (.ZN(I5002A),.A(g1173A));
INV_X1 U_g7550A (.ZN(g7550A),.A(FE_OFN96_g2169A));
INV_X1 U_g2077A (.ZN(g2077A),.A(g219A));
INV_X1 U_g3103A (.ZN(g3103A),.A(g1212A));
INV_X1 U_g7913A (.ZN(g7913A),.A(g7467A));
INV_X1 U_g6109A (.ZN(g6109A),.A(g48A));
INV_X1 U_g6449A (.ZN(g6449A),.A(g5557A));
INV_X1 U_g2273A (.ZN(g2273A),.A(g881A));
INV_X1 U_g7692A (.ZN(g7692A),.A(g2176A));
INV_X1 U_g7497A (.ZN(g7497A),.A(FE_OFN85_g2176A));
INV_X1 U_g2444A (.ZN(g2444A),.A(g876A));
INV_X1 U_g8099A (.ZN(g8099A),.A(g7990A));
INV_X1 U_I9326A (.ZN(I9326A),.A(FE_OFN271_g85A));
INV_X1 U_g6268A (.ZN(g6268A),.A(I9346A));
INV_X1 U_g10676A (.ZN(g10676A),.A(g10570A));
INV_X1 U_g1993A (.ZN(g1993A),.A(g786A));
INV_X1 U_I9383A (.ZN(I9383A),.A(g88A));
INV_X1 U_g8983A (.ZN(g8983A),.A(I14315A));
INV_X1 U_I5254A (.ZN(I5254A),.A(g1700A));
INV_X1 U_I14303A (.ZN(I14303A),.A(g8811A));
INV_X1 U_g2178A (.ZN(g2178A),.A(g45A));
INV_X1 U_I4900A (.ZN(I4900A),.A(g583A));
INV_X1 U_g3060A (.ZN(g3060A),.A(FE_OFN245_g1690A));
INV_X1 U_g4214A (.ZN(g4214A),.A(I5053A));
INV_X1 U_I9346A (.ZN(I9346A),.A(g86A));
INV_X1 U_g2382A (.ZN(g2382A),.A(g599A));
INV_X1 U_g3784A (.ZN(g3784A),.A(FE_OFN254_g461A));
INV_X1 U_I17413A (.ZN(I17413A),.A(g11425A));
INV_X1 U_g7677A (.ZN(g7677A),.A(FE_OFN85_g2176A));
INV_X4 U_g4002A (.ZN(g4002A),.A(FE_OFN155_g3121A));
INV_X1 U_g3479A (.ZN(g3479A),.A(g1101A));
INV_X1 U_g11489A (.ZN(g11489A),.A(I17413A));
INV_X1 U_g6131A (.ZN(g6131A),.A(g5548A));
INV_X1 U_g3390A (.ZN(g3390A),.A(g2045A));
INV_X1 U_g5627A (.ZN(g5627A),.A(FE_OFN132_g3015A));
INV_X1 U_g3501A (.ZN(g3501A),.A(FE_OFN240_g1110A));
INV_X1 U_g8335A (.ZN(g8335A),.A(I13385A));
INV_X1 U_g2095A (.ZN(g2095A),.A(g143A));
INV_X1 U_g2208A (.ZN(g2208A),.A(g84A));
INV_X1 U_g2579A (.ZN(g2579A),.A(g1969A));
INV_X1 U_I14326A (.ZN(I14326A),.A(g8818A));
INV_X1 U_g6283A (.ZN(g6283A),.A(I9311A));
INV_X1 U_g6920A (.ZN(g6920A),.A(I7817A));
INV_X1 U_g8095A (.ZN(g8095A),.A(g7942A));
INV_X1 U_g6718A (.ZN(g6718A),.A(FE_OFN116_g4807A));
INV_X1 U_g2364A (.ZN(g2364A),.A(g611A));
INV_X1 U_g4194A (.ZN(g4194A),.A(I5399A));
INV_X1 U_g2054A (.ZN(g2054A),.A(g1864A));
INV_X1 U_g6261A (.ZN(g6261A),.A(I9265A));
INV_X1 U_g2725A (.ZN(g2725A),.A(g2018A));
INV_X1 U_g5503A (.ZN(g5503A),.A(FE_OFN204_g3664A));
INV_X1 U_g10465A (.ZN(g10465A),.A(I15986A));
INV_X1 U_g1980A (.ZN(g1980A),.A(g646A));
INV_X1 U_g8164A (.ZN(g8164A),.A(g2216A));
INV_X1 U_g8233A (.ZN(g8233A),.A(g2216A));
INV_X1 U_I6220A (.ZN(I6220A),.A(g883A));
INV_X1 U_I4891A (.ZN(I4891A),.A(g582A));
INV_X1 U_I4859A (.ZN(I4859A),.A(g578A));
INV_X1 U_g4212A (.ZN(g4212A),.A(I5044A));
INV_X1 U_I9479A (.ZN(I9479A),.A(g29A));
INV_X1 U_g2297A (.ZN(g2297A),.A(g865A));
INV_X1 U_g7622A (.ZN(g7622A),.A(g7067A));
INV_X1 U_I13400A (.ZN(I13400A),.A(g8236A));
INV_X1 U_g2338A (.ZN(g2338A),.A(g1909A));
INV_X1 U_g7446A (.ZN(g7446A),.A(FE_OFN86_g2176A));
INV_X1 U_g3475A (.ZN(g3475A),.A(g3056A));
INV_X1 U_g4822A (.ZN(g4822A),.A(g3706A));
INV_X1 U_g10437A (.ZN(g10437A),.A(g10333A));
INV_X1 U_g3039A (.ZN(g3039A),.A(g2310A));
INV_X1 U_I6240A (.ZN(I6240A),.A(g878A));
INV_X1 U_I9810A (.ZN(I9810A),.A(g5576A));
INV_X1 U_g2449A (.ZN(g2449A),.A(g790A));
INV_X1 U_I4783A (.ZN(I4783A),.A(g873A));
INV_X1 U_g2604A (.ZN(g2604A),.A(I5525A));
INV_X1 U_I5399A (.ZN(I5399A),.A(g895A));
INV_X1 U_g6165A (.ZN(g6165A),.A(FE_OFN100_g4421A));
INV_X1 U_I5510A (.ZN(I5510A),.A(g588A));
INV_X1 U_I5245A (.ZN(I5245A),.A(g925A));
INV_X1 U_g9505A (.ZN(g9505A),.A(FE_OFN56_g9052A));
INV_X1 U_g2268A (.ZN(g2268A),.A(g654A));
INV_X1 U_g4192A (.ZN(g4192A),.A(I5388A));
INV_X1 U_g3546A (.ZN(g3546A),.A(FE_OFN352_g109A));
INV_X4 U_g9474A (.ZN(g9474A),.A(g9331A));
INV_X1 U_g5222A (.ZN(g5222A),.A(FE_OFN153_g4640A));
INV_X1 U_g2070A (.ZN(g2070A),.A(g213A));
INV_X1 U_g3906A (.ZN(g3906A),.A(FE_OFN364_g3015A));
INV_X1 U_I4866A (.ZN(I4866A),.A(g579A));
INV_X1 U_g6256A (.ZN(g6256A),.A(g2216A));
INV_X1 U_g4176A (.ZN(g4176A),.A(g1989A));
INV_X1 U_g2331A (.ZN(g2331A),.A(g658A));
INV_X1 U_g2406A (.ZN(g2406A),.A(g1365A));
INV_X1 U_I13332A (.ZN(I13332A),.A(g8206A));
INV_X1 U_g6263A (.ZN(g6263A),.A(I9290A));
INV_X1 U_g11239A (.ZN(g11239A),.A(FE_OFN13_g10702A));
INV_X1 U_g2087A (.ZN(g2087A),.A(g225A));
INV_X1 U_g2801A (.ZN(g2801A),.A(g2117A));
INV_X1 U_g3738A (.ZN(g3738A),.A(g3062A));
INV_X1 U_g7512A (.ZN(g7512A),.A(FE_OFN86_g2176A));
INV_X1 U_g9760A (.ZN(g9760A),.A(FE_OFN33_g9454A));
INV_X1 U_g6257A (.ZN(g6257A),.A(g2169A));
INV_X1 U_g4177A (.ZN(g4177A),.A(g1990A));
INV_X1 U_g4206A (.ZN(g4206A),.A(I5579A));
INV_X1 U_g2045A (.ZN(g2045A),.A(g1811A));
INV_X1 U_g8331A (.ZN(g8331A),.A(I13373A));
INV_X1 U_I9276A (.ZN(I9276A),.A(g83A));
INV_X1 U_g8105A (.ZN(g8105A),.A(g7992A));
INV_X1 U_g2169A (.ZN(g2169A),.A(g42A));
INV_X1 U_I5395A (.ZN(I5395A),.A(g892A));
INV_X1 U_g2369A (.ZN(g2369A),.A(g617A));
INV_X1 U_g2602A (.ZN(g2602A),.A(I5497A));
INV_X1 U_g4199A (.ZN(g4199A),.A(I5418A));
INV_X1 U_g2407A (.ZN(g2407A),.A(g197A));
INV_X1 U_g9451A (.ZN(g9451A),.A(I14642A));
INV_X1 U_g5836A (.ZN(g5836A),.A(FE_OFN273_g85A));
INV_X1 U_g4207A (.ZN(g4207A),.A(I5584A));
INV_X1 U_g11083A (.ZN(g11083A),.A(g10788A));
INV_X1 U_g11348A (.ZN(g11348A),.A(g11276A));
INV_X1 U_I5815A (.ZN(I5815A),.A(g794A));
INV_X1 U_g9508A (.ZN(g9508A),.A(g9271A));
INV_X1 U_g2203A (.ZN(g2203A),.A(g677A));
INV_X1 U_g7686A (.ZN(g7686A),.A(FE_OFN85_g2176A));
INV_X1 U_I5497A (.ZN(I5497A),.A(g587A));
INV_X1 U_I13421A (.ZN(I13421A),.A(g8200A));
INV_X1 U_g4215A (.ZN(g4215A),.A(I5060A));
INV_X1 U_g6863A (.ZN(g6863A),.A(g6740A));
INV_X1 U_g2216A (.ZN(g2216A),.A(g41A));
INV_X1 U_g2028A (.ZN(g2028A),.A(g1703A));
INV_X1 U_g4336A (.ZN(g4336A),.A(g4130A));
INV_X1 U_g2564A (.ZN(g2564A),.A(g1814A));
INV_X1 U_g3705A (.ZN(g3705A),.A(FE_OFN308_I6424A));
INV_X1 U_g4065A (.ZN(g4065A),.A(g2794A));
INV_X1 U_g4887A (.ZN(g4887A),.A(I5057A));
INV_X1 U_g2609A (.ZN(g2609A),.A(I4900A));
INV_X1 U_g4934A (.ZN(g4934A),.A(g4243A));
INV_X1 U_g3814A (.ZN(g3814A),.A(g2355A));
INV_X1 U_g8564A (.ZN(g8564A),.A(I7840A));
INV_X1 U_g2571A (.ZN(g2571A),.A(g1822A));
INV_X1 U_g4195A (.ZN(g4195A),.A(I5406A));
INV_X1 U_g1975A (.ZN(g1975A),.A(g622A));
INV_X1 U_g2774A (.ZN(g2774A),.A(FE_OFN225_g2276A));
INV_X1 U_g3967A (.ZN(g3967A),.A(g3247A));
INV_X1 U_I4935A (.ZN(I4935A),.A(g585A));
INV_X1 U_g2396A (.ZN(g2396A),.A(g1389A));
INV_X1 U_g1984A (.ZN(g1984A),.A(g758A));
INV_X1 U_g11539A (.ZN(g11539A),.A(g11519A));
INV_X1 U_g2018A (.ZN(g2018A),.A(g1336A));
INV_X1 U_g2067A (.ZN(g2067A),.A(g108A));
INV_X1 U_I14323A (.ZN(I14323A),.A(g8817A));
INV_X1 U_I14299A (.ZN(I14299A),.A(g8810A));
INV_X1 U_I6277A (.ZN(I6277A),.A(g1206A));
INV_X1 U_I9237A (.ZN(I9237A),.A(g31A));
INV_X1 U_g2381A (.ZN(g2381A),.A(g1368A));
INV_X1 U_g9432A (.ZN(g9432A),.A(g9313A));
INV_X1 U_g8509A (.ZN(g8509A),.A(g8366A));
INV_X1 U_g7905A (.ZN(g7905A),.A(g7450A));
INV_X1 U_g2421A (.ZN(g2421A),.A(g1374A));
INV_X1 U_g4001A (.ZN(g4001A),.A(g3200A));
INV_X1 U_g11515A (.ZN(g11515A),.A(g11490A));
INV_X1 U_g3485A (.ZN(g3485A),.A(g1104A));
INV_X1 U_g2562A (.ZN(g2562A),.A(g1383A));
INV_X1 U_g6697A (.ZN(g6697A),.A(g4807A));
INV_X1 U_g8700A (.ZN(g8700A),.A(g8574A));
INV_X1 U_g2605A (.ZN(g2605A),.A(I4866A));
INV_X1 U_g11206A (.ZN(g11206A),.A(g10629A));
INV_X1 U_I5427A (.ZN(I5427A),.A(g913A));
INV_X1 U_I9769A (.ZN(I9769A),.A(g5287A));
INV_X1 U_g11107A (.ZN(g11107A),.A(FE_OFN7_g10702A));
INV_X1 U_I11360A (.ZN(I11360A),.A(g6351A));
INV_X1 U_g8562A (.ZN(g8562A),.A(I7825A));
INV_X1 U_g9778A (.ZN(g9778A),.A(FE_OFN63_g9474A));
INV_X1 U_g3765A (.ZN(g3765A),.A(g3120A));
INV_X1 U_g4198A (.ZN(g4198A),.A(I5414A));
INV_X1 U_I14330A (.ZN(I14330A),.A(g8819A));
INV_X1 U_g9526A (.ZN(g9526A),.A(g9256A));
INV_X1 U_I15962A (.ZN(I15962A),.A(g10405A));
INV_X1 U_g3069A (.ZN(g3069A),.A(I6277A));
INV_X1 U_I15500A (.ZN(I15500A),.A(g10019A));
INV_X1 U_I5047A (.ZN(I5047A),.A(g1185A));
INV_X1 U_g2074A (.ZN(g2074A),.A(g1377A));
INV_X1 U_I16507A (.ZN(I16507A),.A(g10712A));
INV_X1 U_g6942A (.ZN(g6942A),.A(I7840A));
INV_X1 U_g4211A (.ZN(g4211A),.A(I5041A));
INV_X1 U_g6432A (.ZN(g6432A),.A(FE_OFN219_g5557A));
INV_X1 U_g7908A (.ZN(g7908A),.A(g7454A));
INV_X1 U_g9764A (.ZN(g9764A),.A(FE_OFN59_g9432A));
INV_X1 U_g3291A (.ZN(g3291A),.A(g2161A));
INV_X1 U_g3207A (.ZN(g3207A),.A(g2439A));
INV_X1 U_g2126A (.ZN(g2126A),.A(g12A));
INV_X1 U_I15514A (.ZN(I15514A),.A(g10007A));
INV_X1 U_I15507A (.ZN(I15507A),.A(g10001A));
INV_X1 U_g1964A (.ZN(g1964A),.A(g114A));
INV_X1 U_g10387A (.ZN(g10387A),.A(g10357A));
INV_X1 U_g11163A (.ZN(g11163A),.A(I16717A));
INV_X1 U_g8688A (.ZN(g8688A),.A(g8507A));
INV_X1 U_g8976A (.ZN(g8976A),.A(I14323A));
INV_X1 U_g2608A (.ZN(g2608A),.A(I4891A));
INV_X1 U_g7450A (.ZN(g7450A),.A(FE_OFN87_g2176A));
INV_X1 U_g4200A (.ZN(g4200A),.A(I5424A));
INV_X1 U_g2023A (.ZN(g2023A),.A(g1357A));
INV_X1 U_g7379A (.ZN(g7379A),.A(g6863A));
INV_X1 U_I13427A (.ZN(I13427A),.A(g8241A));
INV_X1 U_I7752A (.ZN(I7752A),.A(g3407A));
INV_X1 U_g4191A (.ZN(g4191A),.A(I5383A));
INV_X1 U_g1989A (.ZN(g1989A),.A(g770A));
INV_X1 U_g3408A (.ZN(g3408A),.A(g3108A));
INV_X1 U_g2451A (.ZN(g2451A),.A(g248A));
INV_X1 U_g8220A (.ZN(g8220A),.A(FE_OFN199_g7697A));
INV_X1 U_g3943A (.ZN(g3943A),.A(g627A));
INV_X1 U_I14295A (.ZN(I14295A),.A(g8806A));
INV_X1 U_g7981A (.ZN(g7981A),.A(g7624A));
INV_X1 U_g6949A (.ZN(g6949A),.A(I7847A));
INV_X1 U_g8977A (.ZN(g8977A),.A(I14295A));
INV_X1 U_g9082A (.ZN(g9082A),.A(FE_OFN76_g8700A));
INV_X1 U_g4811A (.ZN(g4811A),.A(g3661A));
INV_X1 U_g10379A (.ZN(g10379A),.A(I15861A));
INV_X1 U_g7680A (.ZN(g7680A),.A(FE_OFN87_g2176A));
INV_X1 U_g8327A (.ZN(g8327A),.A(g8164A));
INV_X1 U_I13385A (.ZN(I13385A),.A(g8230A));
INV_X1 U_g7744A (.ZN(g7744A),.A(g1962A));
INV_X1 U_g8146A (.ZN(g8146A),.A(FE_OFN330_g7638A));
INV_X1 U_I5057A (.ZN(I5057A),.A(g1961A));
INV_X1 U_I8503A (.ZN(I8503A),.A(FE_OFN184_I7048A));
INV_X1 U_g2034A (.ZN(g2034A),.A(g1766A));
INV_X1 U_g8103A (.ZN(g8103A),.A(g7994A));
INV_X1 U_g2434A (.ZN(g2434A),.A(g1362A));
INV_X1 U_g3913A (.ZN(g3913A),.A(g3121A));
INV_X1 U_g6702A (.ZN(g6702A),.A(FE_OFN117_g4807A));
INV_X1 U_g4880A (.ZN(g4880A),.A(FE_OFN292_g3015A));
INV_X1 U_g8696A (.ZN(g8696A),.A(g8488A));
INV_X1 U_I14309A (.ZN(I14309A),.A(g8813A));
INV_X1 U_g2347A (.ZN(g2347A),.A(g1945A));
INV_X1 U_g6276A (.ZN(g6276A),.A(I9329A));
INV_X1 U_g4243A (.ZN(g4243A),.A(g3524A));
INV_X1 U_I9259A (.ZN(I9259A),.A(g89A));
INV_X1 U_g7574A (.ZN(g7574A),.A(FE_OFN80_g2175A));
INV_X1 U_g8316A (.ZN(g8316A),.A(I13332A));
INV_X1 U_g8565A (.ZN(g8565A),.A(I7847A));
INV_X1 U_g8347A (.ZN(g8347A),.A(I13421A));
INV_X1 U_g1962A (.ZN(g1962A),.A(g27A));
INV_X1 U_g2601A (.ZN(g2601A),.A(I4859A));
INV_X1 U_g4213A (.ZN(g4213A),.A(I5047A));
INV_X1 U_g6277A (.ZN(g6277A),.A(I9349A));
INV_X1 U_g2060A (.ZN(g2060A),.A(g1380A));
INV_X1 U_g6617A (.ZN(g6617A),.A(g6019A));
INV_X1 U_I13338A (.ZN(I13338A),.A(g8210A));
INV_X1 U_I15861A (.ZN(I15861A),.A(g10339A));
INV_X1 U_I5525A (.ZN(I5525A),.A(g589A));
INV_X1 U_g4456A (.ZN(g4456A),.A(FE_OFN234_g2024A));
INV_X1 U_g2479A (.ZN(g2479A),.A(g26A));
INV_X1 U_I16220A (.ZN(I16220A),.A(g10502A));
INV_X1 U_g9814A (.ZN(g9814A),.A(FE_OFN70_g9490A));
INV_X1 U_g3068A (.ZN(g3068A),.A(g2303A));
INV_X1 U_g9773A (.ZN(g9773A),.A(g9474A));
INV_X1 U_g5200A (.ZN(g5200A),.A(g4567A));
INV_X1 U_g4457A (.ZN(g4457A),.A(FE_OFN137_g3829A));
INV_X1 U_g4193A (.ZN(g4193A),.A(I5395A));
INV_X1 U_g10461A (.ZN(g10461A),.A(I15974A));
INV_X1 U_I5020A (.ZN(I5020A),.A(g1176A));
INV_X1 U_g1969A (.ZN(g1969A),.A(g456A));
INV_X1 U_I9293A (.ZN(I9293A),.A(g92A));
INV_X1 U_I9329A (.ZN(I9329A),.A(g94A));
INV_X1 U_g7903A (.ZN(g7903A),.A(g7446A));
INV_X1 U_I9221A (.ZN(I9221A),.A(g30A));
INV_X1 U_g4525A (.ZN(g4525A),.A(FE_OFN229_g3880A));
INV_X1 U_g2475A (.ZN(g2475A),.A(g192A));
INV_X1 U_g1988A (.ZN(g1988A),.A(g766A));
INV_X1 U_g11203A (.ZN(g11203A),.A(FE_OFN20_g10702A));
INV_X1 U_g4158A (.ZN(g4158A),.A(g3304A));
INV_X1 U_g6557A (.ZN(g6557A),.A(FE_OFN217_g5013A));
INV_X1 U_g2603A (.ZN(g2603A),.A(I5510A));
INV_X1 U_I5410A (.ZN(I5410A),.A(g901A));
INV_X1 U_g10459A (.ZN(g10459A),.A(I15968A));
INV_X1 U_I9349A (.ZN(I9349A),.A(g95A));
INV_X1 U_g6955A (.ZN(g6955A),.A(I7852A));
INV_X1 U_I15290A (.ZN(I15290A),.A(g9974A));
INV_X1 U_g6254A (.ZN(g6254A),.A(I9221A));
INV_X1 U_g4174A (.ZN(g4174A),.A(g1987A));
INV_X1 U_g10444A (.ZN(g10444A),.A(g10325A));
INV_X1 U_I14642A (.ZN(I14642A),.A(g9088A));
INV_X1 U_g4180A (.ZN(g4180A),.A(g1993A));
INV_X1 U_g7917A (.ZN(g7917A),.A(g7497A));
INV_X1 U_g2986A (.ZN(g2986A),.A(I6220A));
INV_X1 U_g9473A (.ZN(g9473A),.A(g9082A));
INV_X1 U_g1965A (.ZN(g1965A),.A(g119A));
INV_X1 U_g11547A (.ZN(g11547A),.A(FE_OFN27_g11519A));
INV_X1 U_g2503A (.ZN(g2503A),.A(g1872A));
INV_X1 U_I9352A (.ZN(I9352A),.A(g28A));
INV_X1 U_I9717A (.ZN(I9717A),.A(FE_OFN97_I8869A));
INV_X1 U_g2224A (.ZN(g2224A),.A(g695A));
INV_X1 U_g7454A (.ZN(g7454A),.A(g2176A));
INV_X1 U_g4204A (.ZN(g4204A),.A(I5445A));
INV_X1 U_g8561A (.ZN(g8561A),.A(I7817A));
INV_X1 U_g8986A (.ZN(g8986A),.A(I14330A));
INV_X1 U_I15956A (.ZN(I15956A),.A(g10402A));
INV_X1 U_I15980A (.ZN(I15980A),.A(g10414A));
AND2_X1 U_g11103A (.ZN(g11103A),.A2(g10937A),.A1(g2250A));
AND2_X1 U_g9900A (.ZN(g9900A),.A2(g8327A),.A1(g9088A));
AND2_X1 U_g11095A (.ZN(g11095A),.A2(FE_OFN4_g10950A),.A1(g845A));
AND2_X2 U_g3880A (.ZN(g3880A),.A2(g2023A),.A1(FE_OFN235_g2024A));
AND2_X1 U_g4973A (.ZN(g4973A),.A2(g4467A),.A1(g1645A));
AND2_X1 U_g7389A (.ZN(g7389A),.A2(FE_OFN226_g3880A),.A1(g5852A));
AND2_X1 U_g7888A (.ZN(g7888A),.A2(FE_OFN334_g7045A),.A1(g7465A));
AND2_X1 U_g4969A (.ZN(g4969A),.A2(g4457A),.A1(g1642A));
AND2_X1 U_g8224A (.ZN(g8224A),.A2(g7949A),.A1(g1882A));
AND2_X1 U_g2892A (.ZN(g2892A),.A2(g1976A),.A1(g1980A));
AND2_X1 U_g5686A (.ZN(g5686A),.A2(FE_OFN365_g5361A),.A1(g158A));
AND2_X1 U_g10308A (.ZN(g10308A),.A2(g9082A),.A1(g10013A));
AND2_X1 U_g4123A (.ZN(g4123A),.A2(g2424A),.A1(g1781A));
AND2_X1 U_g8120A (.ZN(g8120A),.A2(g7949A),.A1(g1909A));
AND2_X1 U_g6788A (.ZN(g6788A),.A2(FE_OFN320_g5361A),.A1(g287A));
AND2_X1 U_g5598A (.ZN(g5598A),.A2(g4824A),.A1(g778A));
AND2_X1 U_g9694A (.ZN(g9694A),.A2(FE_OFN59_g9432A),.A1(g278A));
AND2_X1 U_g10495A (.ZN(g10495A),.A2(FE_OFN234_g2024A),.A1(g10431A));
AND2_X1 U_g2945A (.ZN(g2945A),.A2(g1684A),.A1(FE_OFN241_g1690A));
AND2_X1 U_g11190A (.ZN(g11190A),.A2(g10927A),.A1(g4752A));
AND2_X1 U_g8789A (.ZN(g8789A),.A2(FE_OFN331_g8696A),.A1(g8639A));
AND2_X1 U_g9852A (.ZN(g9852A),.A2(g9563A),.A1(g9728A));
AND2_X1 U_g5625A (.ZN(g5625A),.A2(g5627A),.A1(g1053A));
AND2_X1 U_g4875A (.ZN(g4875A),.A2(g4673A),.A1(g995A));
AND2_X1 U_g9701A (.ZN(g9701A),.A2(g9474A),.A1(g1574A));
AND2_X1 U_g7138A (.ZN(g7138A),.A2(g6718A),.A1(g5201A));
AND2_X1 U_g10752A (.ZN(g10752A),.A2(FE_OFN103_g3586A),.A1(g10599A));
AND2_X1 U_g11211A (.ZN(g11211A),.A2(g5503A),.A1(g11058A));
AND2_X1 U_g11024A (.ZN(g11024A),.A2(g10702A),.A1(g435A));
AND2_X1 U_g8547A (.ZN(g8547A),.A2(FE_OFN211_g7246A),.A1(g8307A));
AND2_X1 U_g10669A (.ZN(g10669A),.A2(g9473A),.A1(g10408A));
AND2_X1 U_g7707A (.ZN(g7707A),.A2(FE_OFN191_g6488A),.A1(g691A));
AND2_X1 U_g4884A (.ZN(g4884A),.A2(g1845A),.A1(g3813A));
AND2_X1 U_g4839A (.ZN(g4839A),.A2(g2355A),.A1(g225A));
AND2_X1 U_g9870A (.ZN(g9870A),.A2(g9802A),.A1(g1561A));
AND2_X1 U_g6640A (.ZN(g6640A),.A2(g5808A),.A1(g86A));
AND2_X1 U_g9650A (.ZN(g9650A),.A2(FE_OFN40_g9240A),.A1(g986A));
AND2_X1 U_g5687A (.ZN(g5687A),.A2(FE_OFN365_g5361A),.A1(g139A));
AND2_X1 U_g7957A (.ZN(g7957A),.A2(g7527A),.A1(g79A));
AND2_X1 U_g3512A (.ZN(g3512A),.A2(g1845A),.A1(g2050A));
AND2_X1 U_g8244A (.ZN(g8244A),.A2(FE_OFN310_g4336A),.A1(g7054A));
AND2_X1 U_g7449A (.ZN(g7449A),.A2(FE_OFN221_g3440A),.A1(g6548A));
AND2_X1 U_g4235A (.ZN(g4235A),.A2(FE_OFN347_g3914A),.A1(g1011A));
AND2_X1 U_g4343A (.ZN(g4343A),.A2(FE_OFN287_g3586A),.A1(g345A));
AND2_X1 U_g11296A (.ZN(g11296A),.A2(g11239A),.A1(g4561A));
AND2_X1 U_g9594A (.ZN(g9594A),.A2(g9292A),.A1(g1A));
AND2_X1 U_g6829A (.ZN(g6829A),.A2(FE_OFN179_g5354A),.A1(g213A));
AND2_X1 U_g4334A (.ZN(g4334A),.A2(FE_OFN351_g3913A),.A1(g1160A));
AND2_X1 U_g9943A (.ZN(g9943A),.A2(FE_OFN67_g9367A),.A1(g9923A));
AND2_X1 U_g5525A (.ZN(g5525A),.A2(g4292A),.A1(g1721A));
AND2_X1 U_g4548A (.ZN(g4548A),.A2(g4002A),.A1(g440A));
AND3_X1 U_g8876A (.ZN(g8876A),.A3(FE_OFN73_g8858A),.A2(FE_OFN93_g2216A),.A1(g8105A));
AND2_X1 U_g6733A (.ZN(g6733A),.A2(FE_OFN322_g4449A),.A1(g4488A));
AND2_X1 U_g4804A (.ZN(g4804A),.A2(g4010A),.A1(g476A));
AND2_X1 U_g10705A (.ZN(g10705A),.A2(FE_OFN131_g3015A),.A1(g10564A));
AND2_X1 U_g9934A (.ZN(g9934A),.A2(g9624A),.A1(g9913A));
AND2_X1 U_g6225A (.ZN(g6225A),.A2(g5613A),.A1(g566A));
AND2_X1 U_g6324A (.ZN(g6324A),.A2(FE_OFN116_g4807A),.A1(g1240A));
AND2_X1 U_g10686A (.ZN(g10686A),.A2(FE_OFN136_g3863A),.A1(g10385A));
AND2_X1 U_g6540A (.ZN(g6540A),.A2(g6081A),.A1(g1223A));
AND2_X1 U_g8663A (.ZN(g8663A),.A2(FE_OFN292_g3015A),.A1(g8270A));
AND2_X1 U_g11581A (.ZN(g11581A),.A2(g11539A),.A1(g1308A));
AND2_X1 U_g6206A (.ZN(g6206A),.A2(g5613A),.A1(g560A));
AND2_X1 U_g4518A (.ZN(g4518A),.A2(g4002A),.A1(g452A));
AND2_X1 U_g3989A (.ZN(g3989A),.A2(FE_OFN359_g18A),.A1(g248A));
AND2_X1 U_g7730A (.ZN(g7730A),.A2(g2347A),.A1(g7260A));
AND2_X1 U_g5174A (.ZN(g5174A),.A2(FE_OFN303_g4678A),.A1(g1235A));
AND2_X1 U_g7504A (.ZN(g7504A),.A2(g67A),.A1(FE_OFN86_g2176A));
AND2_X1 U_g7185A (.ZN(g7185A),.A2(FE_OFN213_g6003A),.A1(g1887A));
AND2_X1 U_g2563A (.ZN(g2563A),.A2(I5690A),.A1(I5689A));
AND2_X1 U_g7881A (.ZN(g7881A),.A2(FE_OFN366_g3521A),.A1(g5295A));
AND2_X1 U_g11070A (.ZN(g11070A),.A2(g10788A),.A1(g2008A));
AND2_X1 U_g9859A (.ZN(g9859A),.A2(g9579A),.A1(g9736A));
AND3_X1 U_g8877A (.ZN(g8877A),.A3(FE_OFN73_g8858A),.A2(FE_OFN92_g2216A),.A1(g8103A));
AND2_X1 U_g11590A (.ZN(g11590A),.A2(g11561A),.A1(g2274A));
AND2_X1 U_g6199A (.ZN(g6199A),.A2(FE_OFN289_g4679A),.A1(g557A));
AND2_X1 U_g9266A (.ZN(g9266A),.A2(FE_OFN325_g18A),.A1(g8932A));
AND2_X1 U_g5545A (.ZN(g5545A),.A2(g4292A),.A1(g1730A));
AND2_X1 U_g5180A (.ZN(g5180A),.A2(g810A),.A1(g814A));
AND2_X1 U_g5591A (.ZN(g5591A),.A2(FE_OFN367_g3521A),.A1(g1615A));
AND2_X1 U_g8556A (.ZN(g8556A),.A2(FE_OFN189_g7638A),.A1(g8412A));
AND2_X1 U_g11094A (.ZN(g11094A),.A2(g10883A),.A1(g374A));
AND2_X1 U_g5853A (.ZN(g5853A),.A2(g1927A),.A1(g5044A));
AND2_X1 U_g6245A (.ZN(g6245A),.A2(FE_OFN289_g4679A),.A1(g575A));
AND2_X1 U_g4360A (.ZN(g4360A),.A2(g3523A),.A1(g1861A));
AND3_X1 U_g8930A (.ZN(g8930A),.A3(g8828A),.A2(FE_OFN95_g2216A),.A1(g8100A));
AND2_X1 U_g5507A (.ZN(g5507A),.A2(FE_OFN357_g3521A),.A1(g563A));
AND2_X1 U_g11150A (.ZN(g11150A),.A2(g10788A),.A1(g3087A));
AND2_X1 U_g8464A (.ZN(g8464A),.A2(FE_OFN210_g7246A),.A1(g8302A));
AND2_X1 U_g9692A (.ZN(g9692A),.A2(FE_OFN59_g9432A),.A1(g272A));
AND2_X1 U_g4996A (.ZN(g4996A),.A2(FE_OFN146_g4682A),.A1(g1428A));
AND2_X1 U_g7131A (.ZN(g7131A),.A2(g6702A),.A1(g5174A));
AND2_X1 U_g11019A (.ZN(g11019A),.A2(FE_OFN7_g10702A),.A1(g421A));
AND2_X1 U_g9960A (.ZN(g9960A),.A2(FE_OFN280_g9536A),.A1(g9951A));
AND2_X1 U_g11196A (.ZN(g11196A),.A2(FE_OFN15_g10702A),.A1(g4770A));
AND2_X1 U_g11018A (.ZN(g11018A),.A2(FE_OFN7_g10702A),.A1(g6485A));
AND2_X1 U_g6819A (.ZN(g6819A),.A2(FE_OFN179_g5354A),.A1(g243A));
AND2_X1 U_g10595A (.ZN(g10595A),.A2(FE_OFN369_g4525A),.A1(g10550A));
AND2_X1 U_g10494A (.ZN(g10494A),.A2(g2024A),.A1(g10433A));
AND2_X1 U_g10623A (.ZN(g10623A),.A2(FE_OFN370_g4525A),.A1(g10544A));
AND2_X1 U_g4878A (.ZN(g4878A),.A2(g3523A),.A1(g1868A));
AND2_X1 U_g5204A (.ZN(g5204A),.A2(g2126A),.A1(g4838A));
AND2_X1 U_g8844A (.ZN(g8844A),.A2(g8709A),.A1(g8609A));
AND2_X1 U_g6701A (.ZN(g6701A),.A2(g4381A),.A1(g6185A));
AND2_X1 U_g10782A (.ZN(g10782A),.A2(g4467A),.A1(g10725A));
AND2_X1 U_g5100A (.ZN(g5100A),.A2(g4608A),.A1(g1791A));
AND2_X1 U_g4882A (.ZN(g4882A),.A2(FE_OFN293_g3015A),.A1(g1089A));
AND2_X1 U_g8731A (.ZN(g8731A),.A2(g7918A),.A1(g8236A));
AND2_X1 U_g6215A (.ZN(g6215A),.A2(g5128A),.A1(g1504A));
AND2_X1 U_g6886A (.ZN(g6886A),.A2(FE_OFN213_g6003A),.A1(g1932A));
AND2_X4 U_g3586A (.ZN(g3586A),.A2(I6260A),.A1(g1703A));
AND2_X1 U_g8557A (.ZN(g8557A),.A2(g7638A),.A1(g8415A));
AND3_X1 U_g8966A (.ZN(g8966A),.A3(g8849A),.A2(FE_OFN93_g2216A),.A1(g8081A));
AND2_X1 U_g8071A (.ZN(g8071A),.A2(FE_OFN199_g7697A),.A1(g691A));
AND2_X1 U_g11597A (.ZN(g11597A),.A2(FE_OFN99_g4421A),.A1(g11549A));
AND2_X1 U_g9828A (.ZN(g9828A),.A2(g9785A),.A1(g9722A));
AND2_X1 U_g2918A (.ZN(g2918A),.A2(g1672A),.A1(FE_OFN241_g1690A));
AND2_X1 U_g9830A (.ZN(g9830A),.A2(FE_OFN34_g9785A),.A1(g9725A));
AND3_X1 U_g8955A (.ZN(g8955A),.A3(g8828A),.A2(FE_OFN95_g2216A),.A1(g8110A));
AND2_X1 U_g9592A (.ZN(g9592A),.A2(g9292A),.A1(g4A));
AND2_X1 U_g5123A (.ZN(g5123A),.A2(g3906A),.A1(g1618A));
AND2_X1 U_g7059A (.ZN(g7059A),.A2(g6354A),.A1(g6078A));
AND2_X1 U_g8254A (.ZN(g8254A),.A2(g7907A),.A1(g936A));
AND2_X1 U_g7459A (.ZN(g7459A),.A2(g55A),.A1(FE_OFN86_g2176A));
AND2_X1 U_g11102A (.ZN(g11102A),.A2(FE_OFN3_g10950A),.A1(g861A));
AND2_X1 U_g7718A (.ZN(g7718A),.A2(FE_OFN191_g6488A),.A1(g709A));
AND2_X1 U_g7535A (.ZN(g7535A),.A2(g49A),.A1(FE_OFN86_g2176A));
AND2_X1 U_g9703A (.ZN(g9703A),.A2(g9474A),.A1(g1577A));
AND2_X1 U_g5528A (.ZN(g5528A),.A2(FE_OFN357_g3521A),.A1(g569A));
AND2_X1 U_g9932A (.ZN(g9932A),.A2(g9624A),.A1(g9911A));
AND2_X1 U_g5530A (.ZN(g5530A),.A2(FE_OFN290_g4880A),.A1(g1636A));
AND2_X1 U_g3506A (.ZN(g3506A),.A2(g2760A),.A1(g986A));
AND2_X1 U_g8769A (.ZN(g8769A),.A2(FE_OFN304_g5151A),.A1(g8629A));
AND2_X1 U_g6887A (.ZN(g6887A),.A2(g6557A),.A1(g6187A));
AND2_X1 U_g6228A (.ZN(g6228A),.A2(g713A),.A1(g5605A));
AND2_X1 U_g6322A (.ZN(g6322A),.A2(FE_OFN116_g4807A),.A1(g1275A));
AND2_X1 U_g3111A (.ZN(g3111A),.A2(I6338A),.A1(I6337A));
AND3_X1 U_g8967A (.ZN(g8967A),.A3(g8849A),.A2(FE_OFN281_g2216A),.A1(g8085A));
AND2_X1 U_g5010A (.ZN(g5010A),.A2(FE_OFN153_g4640A),.A1(g1458A));
AND2_X1 U_g3275A (.ZN(g3275A),.A2(FE_OFN266_g18A),.A1(g115A));
AND2_X1 U_g10809A (.ZN(g10809A),.A2(g10702A),.A1(g4811A));
AND2_X1 U_g2895A (.ZN(g2895A),.A2(g1678A),.A1(FE_OFN336_g1690A));
AND2_X1 U_g7721A (.ZN(g7721A),.A2(g6488A),.A1(g736A));
AND2_X1 U_g9866A (.ZN(g9866A),.A2(g9802A),.A1(g1549A));
AND2_X1 U_g9716A (.ZN(g9716A),.A2(FE_OFN70_g9490A),.A1(g1534A));
AND2_X1 U_g10808A (.ZN(g10808A),.A2(FE_OFN137_g3829A),.A1(g10744A));
AND2_X1 U_g3374A (.ZN(g3374A),.A2(g3047A),.A1(g1231A));
AND2_X1 U_g4492A (.ZN(g4492A),.A2(g3685A),.A1(FE_OFN253_g1786A));
AND2_X1 U_g8822A (.ZN(g8822A),.A2(FE_OFN328_g8709A),.A1(g8614A));
AND2_X1 U_g10560A (.ZN(g10560A),.A2(FE_OFN369_g4525A),.A1(g10369A));
AND3_X1 U_g11456A (.ZN(g11456A),.A3(g11348A),.A2(g2801A),.A1(g3765A));
AND2_X1 U_g9848A (.ZN(g9848A),.A2(g9579A),.A1(g9724A));
AND2_X1 U_g4714A (.ZN(g4714A),.A2(g3943A),.A1(g646A));
AND2_X1 U_g6550A (.ZN(g6550A),.A2(g6081A),.A1(g1231A));
AND2_X1 U_g5172A (.ZN(g5172A),.A2(g818A),.A1(g822A));
AND2_X1 U_g10642A (.ZN(g10642A),.A2(g3829A),.A1(g10385A));
AND2_X1 U_g3284A (.ZN(g3284A),.A2(g677A),.A1(g2531A));
AND2_X1 U_g9699A (.ZN(g9699A),.A2(FE_OFN59_g9432A),.A1(g284A));
AND2_X1 U_g9855A (.ZN(g9855A),.A2(g9764A),.A1(g302A));
AND2_X1 U_g5618A (.ZN(g5618A),.A2(FE_OFN367_g3521A),.A1(g1630A));
AND2_X1 U_g6891A (.ZN(g6891A),.A2(g6003A),.A1(g1950A));
AND2_X1 U_g7940A (.ZN(g7940A),.A2(FE_OFN292_g3015A),.A1(g5319A));
AND2_X1 U_g11085A (.ZN(g11085A),.A2(g10927A),.A1(g312A));
AND2_X1 U_g4736A (.ZN(g4736A),.A2(FE_OFN300_g4002A),.A1(g396A));
AND2_X1 U_g4968A (.ZN(g4968A),.A2(FE_OFN146_g4682A),.A1(g1432A));
AND2_X1 U_g8837A (.ZN(g8837A),.A2(FE_OFN331_g8696A),.A1(g8646A));
AND2_X1 U_g9644A (.ZN(g9644A),.A2(FE_OFN45_g9125A),.A1(g1182A));
AND2_X1 U_g5804A (.ZN(g5804A),.A2(g5261A),.A1(g1546A));
AND2_X1 U_g8462A (.ZN(g8462A),.A2(FE_OFN211_g7246A),.A1(g8300A));
AND4_X1 U_I6330A (.ZN(I6330A),.A4(g2570A),.A3(g2562A),.A2(g2556A),.A1(g2549A));
AND2_X1 U_g11156A (.ZN(g11156A),.A2(FE_OFN278_g10927A),.A1(g333A));
AND2_X1 U_g6342A (.ZN(g6342A),.A2(FE_OFN319_g5361A),.A1(g293A));
AND2_X1 U_g9867A (.ZN(g9867A),.A2(g9802A),.A1(g1552A));
AND2_X1 U_g9717A (.ZN(g9717A),.A2(FE_OFN70_g9490A),.A1(g1537A));
AND2_X1 U_g4871A (.ZN(g4871A),.A2(g3523A),.A1(g1864A));
AND2_X1 U_g10454A (.ZN(g10454A),.A2(FE_OFN235_g2024A),.A1(g10435A));
AND2_X1 U_g4722A (.ZN(g4722A),.A2(FE_OFN300_g4002A),.A1(g426A));
AND2_X1 U_g7741A (.ZN(g7741A),.A2(g3880A),.A1(g5824A));
AND2_X1 U_g4500A (.ZN(g4500A),.A2(FE_OFN291_g4880A),.A1(g1357A));
AND2_X1 U_g9386A (.ZN(g9386A),.A2(FE_OFN47_g9151A),.A1(g1327A));
AND2_X1 U_g8842A (.ZN(g8842A),.A2(FE_OFN328_g8709A),.A1(g8607A));
AND2_X1 U_g9599A (.ZN(g9599A),.A2(FE_OFN71_g9292A),.A1(g8A));
AND2_X4 U_g9274A (.ZN(g9274A),.A2(FE_OFN275_g48A),.A1(g8974A));
AND2_X1 U_g5518A (.ZN(g5518A),.A2(FE_OFN357_g3521A),.A1(g566A));
AND2_X1 U_g9614A (.ZN(g9614A),.A2(FE_OFN51_g9111A),.A1(g1197A));
AND2_X1 U_g4838A (.ZN(g4838A),.A2(g4122A),.A1(g3275A));
AND2_X4 U_g9125A (.ZN(g9125A),.A2(FE_OFN276_g48A),.A1(g8966A));
AND2_X1 U_g7217A (.ZN(g7217A),.A2(g6432A),.A1(g4610A));
AND2_X1 U_g11557A (.ZN(g11557A),.A2(g11519A),.A1(g1791A));
AND2_X1 U_g2911A (.ZN(g2911A),.A2(g1675A),.A1(FE_OFN336_g1690A));
AND2_X1 U_g11210A (.ZN(g11210A),.A2(FE_OFN204_g3664A),.A1(g10886A));
AND2_X1 U_g7466A (.ZN(g7466A),.A2(g58A),.A1(g2176A));
AND2_X1 U_g9939A (.ZN(g9939A),.A2(FE_OFN67_g9367A),.A1(g9918A));
AND2_X1 U_g11279A (.ZN(g11279A),.A2(g11203A),.A1(g4784A));
AND3_X1 U_g10518A (.ZN(g10518A),.A3(I16145A),.A2(g10440A),.A1(g10513A));
AND2_X1 U_g4477A (.ZN(g4477A),.A2(g3913A),.A1(g1129A));
AND2_X1 U_g7055A (.ZN(g7055A),.A2(g6586A),.A1(g5004A));
AND2_X1 U_g5264A (.ZN(g5264A),.A2(g4776A),.A1(g1095A));
AND2_X1 U_g6329A (.ZN(g6329A),.A2(FE_OFN115_g4807A),.A1(g1265A));
AND2_X1 U_g6828A (.ZN(g6828A),.A2(FE_OFN179_g5354A),.A1(g1377A));
AND2_X1 U_g8176A (.ZN(g8176A),.A2(FE_OFN89_I11360A),.A1(g40A));
AND2_X1 U_g6830A (.ZN(g6830A),.A2(FE_OFN179_g5354A),.A1(g1380A));
AND2_X1 U_g8005A (.ZN(g8005A),.A2(FE_OFN334_g7045A),.A1(g7510A));
AND2_X1 U_g4099A (.ZN(g4099A),.A2(g3281A),.A1(g770A));
AND2_X1 U_g11601A (.ZN(g11601A),.A2(g11575A),.A1(g1351A));
AND2_X1 U_g11187A (.ZN(g11187A),.A2(FE_OFN10_g10702A),.A1(g4727A));
AND2_X1 U_g6746A (.ZN(g6746A),.A2(FE_OFN218_g5557A),.A1(g6228A));
AND2_X1 U_g6221A (.ZN(g6221A),.A2(g5598A),.A1(g782A));
AND2_X1 U_g8765A (.ZN(g8765A),.A2(FE_OFN304_g5151A),.A1(g8630A));
AND2_X1 U_g9622A (.ZN(g9622A),.A2(FE_OFN51_g9111A),.A1(g1200A));
AND2_X1 U_g11143A (.ZN(g11143A),.A2(g4567A),.A1(g10923A));
AND2_X1 U_g9904A (.ZN(g9904A),.A2(g9676A),.A1(g9886A));
AND2_X1 U_g8733A (.ZN(g8733A),.A2(g7920A),.A1(g8241A));
AND3_X1 U_g8974A (.ZN(g8974A),.A3(FE_OFN73_g8858A),.A2(FE_OFN93_g2216A),.A1(g8094A));
AND2_X1 U_g6624A (.ZN(g6624A),.A2(FE_OFN282_g6165A),.A1(g348A));
AND2_X1 U_g11169A (.ZN(g11169A),.A2(FE_OFN8_g10702A),.A1(g530A));
AND2_X1 U_g8073A (.ZN(g8073A),.A2(FE_OFN199_g7697A),.A1(g709A));
AND2_X1 U_g9841A (.ZN(g9841A),.A2(g9512A),.A1(g9706A));
AND2_X1 U_g5882A (.ZN(g5882A),.A2(FE_OFN141_g3829A),.A1(g5592A));
AND2_X1 U_g8796A (.ZN(g8796A),.A2(FE_OFN331_g8696A),.A1(g8645A));
AND2_X1 U_g11168A (.ZN(g11168A),.A2(FE_OFN7_g10702A),.A1(g534A));
AND2_X1 U_g4269A (.ZN(g4269A),.A2(FE_OFN347_g3914A),.A1(g1015A));
AND2_X1 U_g5271A (.ZN(g5271A),.A2(FE_OFN335_g4737A),.A1(g727A));
AND2_X1 U_g10348A (.ZN(g10348A),.A2(g3705A),.A1(I15500A));
AND2_X1 U_g5611A (.ZN(g5611A),.A2(g4880A),.A1(g1047A));
AND2_X1 U_g8069A (.ZN(g8069A),.A2(FE_OFN198_g7697A),.A1(g673A));
AND2_X1 U_g9695A (.ZN(g9695A),.A2(g9474A),.A1(g1567A));
AND2_X1 U_g10304A (.ZN(g10304A),.A2(g9291A),.A1(g10001A));
AND2_X1 U_g8469A (.ZN(g8469A),.A2(FE_OFN211_g7246A),.A1(g8305A));
AND2_X1 U_g4712A (.ZN(g4712A),.A2(FE_OFN297_g3015A),.A1(g1071A));
AND2_X1 U_g6576A (.ZN(g6576A),.A2(g5503A),.A1(g5762A));
AND2_X1 U_g10622A (.ZN(g10622A),.A2(FE_OFN369_g4525A),.A1(g10496A));
AND2_X1 U_g11015A (.ZN(g11015A),.A2(FE_OFN18_g10702A),.A1(g5217A));
AND2_X1 U_g5674A (.ZN(g5674A),.A2(FE_OFN365_g5361A),.A1(g148A));
AND2_X1 U_g9359A (.ZN(g9359A),.A2(FE_OFN52_g9173A),.A1(g1308A));
AND2_X2 U_g9223A (.ZN(g9223A),.A2(g8960A),.A1(FE_OFN277_g48A));
AND2_X1 U_g11556A (.ZN(g11556A),.A2(g11519A),.A1(g1786A));
AND2_X1 U_g9858A (.ZN(g9858A),.A2(g9778A),.A1(g1595A));
AND2_X1 U_g5541A (.ZN(g5541A),.A2(g3521A),.A1(g575A));
AND2_X1 U_g4534A (.ZN(g4534A),.A2(FE_OFN344_g3586A),.A1(g363A));
AND2_X1 U_g6198A (.ZN(g6198A),.A2(g5128A),.A1(g1499A));
AND2_X1 U_g6747A (.ZN(g6747A),.A2(g5897A),.A1(g2214A));
AND2_X1 U_g6699A (.ZN(g6699A),.A2(FE_OFN111_g3914A),.A1(g6177A));
AND2_X1 U_g6855A (.ZN(g6855A),.A2(g6392A),.A1(g1964A));
AND2_X1 U_g3804A (.ZN(g3804A),.A2(g2203A),.A1(g3098A));
AND2_X1 U_g5680A (.ZN(g5680A),.A2(FE_OFN164_g5361A),.A1(g153A));
AND2_X1 U_g9642A (.ZN(g9642A),.A2(FE_OFN40_g9240A),.A1(g981A));
AND2_X1 U_g5744A (.ZN(g5744A),.A2(FE_OFN321_g5261A),.A1(g1528A));
AND2_X1 U_g10333A (.ZN(g10333A),.A2(FE_OFN267_g109A),.A1(I15500A));
AND2_X1 U_g8399A (.ZN(g8399A),.A2(g8220A),.A1(g5266A));
AND2_X1 U_g9447A (.ZN(g9447A),.A2(FE_OFN49_g9030A),.A1(g1762A));
AND2_X1 U_g4903A (.ZN(g4903A),.A2(g4243A),.A1(g1849A));
AND2_X1 U_g11178A (.ZN(g11178A),.A2(FE_OFN13_g10702A),.A1(g516A));
AND2_X1 U_g8510A (.ZN(g8510A),.A2(FE_OFN330_g7638A),.A1(g8414A));
AND2_X1 U_g8245A (.ZN(g8245A),.A2(FE_OFN322_g4449A),.A1(g7062A));
AND2_X1 U_g6319A (.ZN(g6319A),.A2(FE_OFN118_g4807A),.A1(g1296A));
AND2_X1 U_g11186A (.ZN(g11186A),.A2(FE_OFN10_g10702A),.A1(g4722A));
AND2_X1 U_g2951A (.ZN(g2951A),.A2(g1681A),.A1(FE_OFN241_g1690A));
AND2_X1 U_g6352A (.ZN(g6352A),.A2(FE_OFN319_g5361A),.A1(g278A));
AND2_X1 U_g9595A (.ZN(g9595A),.A2(FE_OFN42_g9205A),.A1(g901A));
AND2_X1 U_g4831A (.ZN(g4831A),.A2(g4109A),.A1(g810A));
AND2_X1 U_g5492A (.ZN(g5492A),.A2(g4263A),.A1(g1654A));
AND2_X1 U_g9272A (.ZN(g9272A),.A2(FE_OFN266_g18A),.A1(g8934A));
AND2_X1 U_g10312A (.ZN(g10312A),.A2(g9082A),.A1(g10019A));
AND2_X1 U_g6186A (.ZN(g6186A),.A2(FE_OFN291_g4880A),.A1(g546A));
AND2_X1 U_g9612A (.ZN(g9612A),.A2(FE_OFN40_g9240A),.A1(g2652A));
AND2_X1 U_g9417A (.ZN(g9417A),.A2(FE_OFN56_g9052A),.A1(g1738A));
AND2_X1 U_g9935A (.ZN(g9935A),.A2(FE_OFN60_g9624A),.A1(g9914A));
AND2_X1 U_g10745A (.ZN(g10745A),.A2(FE_OFN102_g3586A),.A1(g10658A));
AND2_X1 U_g11216A (.ZN(g11216A),.A2(FE_OFN279_g11157A),.A1(g956A));
AND2_X1 U_g9328A (.ZN(g9328A),.A2(FE_OFN275_g48A),.A1(g8971A));
AND2_X1 U_g11587A (.ZN(g11587A),.A2(g11539A),.A1(g1327A));
AND2_X1 U_g6821A (.ZN(g6821A),.A2(FE_OFN178_g5354A),.A1(g237A));
AND2_X1 U_g6325A (.ZN(g6325A),.A2(FE_OFN116_g4807A),.A1(g1245A));
AND2_X1 U_g4560A (.ZN(g4560A),.A2(g4002A),.A1(g431A));
AND2_X1 U_g7368A (.ZN(g7368A),.A2(g3880A),.A1(g5842A));
AND2_X1 U_g6083A (.ZN(g6083A),.A2(g4273A),.A1(g552A));
AND2_X1 U_g6544A (.ZN(g6544A),.A2(g6081A),.A1(g1227A));
AND2_X1 U_g5476A (.ZN(g5476A),.A2(g4673A),.A1(g1615A));
AND2_X1 U_g7743A (.ZN(g7743A),.A2(FE_OFN226_g3880A),.A1(g5838A));
AND2_X1 U_g4869A (.ZN(g4869A),.A2(FE_OFN132_g3015A),.A1(g1083A));
AND2_X1 U_g5722A (.ZN(g5722A),.A2(FE_OFN315_g5117A),.A1(g1598A));
AND2_X1 U_g6790A (.ZN(g6790A),.A2(FE_OFN346_g4381A),.A1(g5813A));
AND2_X1 U_g8408A (.ZN(g8408A),.A2(g8146A),.A1(g704A));
AND2_X1 U_g10761A (.ZN(g10761A),.A2(g10558A),.A1(g10559A));
AND2_X1 U_g7734A (.ZN(g7734A),.A2(FE_OFN226_g3880A),.A1(g5810A));
AND2_X1 U_g8136A (.ZN(g8136A),.A2(g7045A),.A1(g7926A));
AND2_X1 U_g6187A (.ZN(g6187A),.A2(g2340A),.A1(g5569A));
AND2_X1 U_g4752A (.ZN(g4752A),.A2(FE_OFN300_g4002A),.A1(g401A));
AND2_X1 U_g9902A (.ZN(g9902A),.A2(FE_OFN69_g9392A),.A1(g9720A));
AND2_X1 U_g8768A (.ZN(g8768A),.A2(FE_OFN304_g5151A),.A1(g8623A));
AND2_X1 U_g5500A (.ZN(g5500A),.A2(g4281A),.A1(g1657A));
AND2_X1 U_g2496A (.ZN(g2496A),.A2(g369A),.A1(g374A));
AND2_X1 U_g6756A (.ZN(g6756A),.A2(g5877A),.A1(g3010A));
AND3_X1 U_g8972A (.ZN(g8972A),.A3(FE_OFN73_g8858A),.A2(FE_OFN281_g2216A),.A1(g8085A));
AND2_X1 U_g6622A (.ZN(g6622A),.A2(g6165A),.A1(g336A));
AND2_X1 U_g11639A (.ZN(g11639A),.A2(g7897A),.A1(g11612A));
AND2_X1 U_g9366A (.ZN(g9366A),.A2(FE_OFN53_g9173A),.A1(g1311A));
AND2_X1 U_g11230A (.ZN(g11230A),.A2(g11060A),.A1(g471A));
AND2_X1 U_g10328A (.ZN(g10328A),.A2(FE_OFN269_g109A),.A1(I15507A));
AND2_X1 U_g5024A (.ZN(g5024A),.A2(FE_OFN303_g4678A),.A1(g1284A));
AND2_X1 U_g4364A (.ZN(g4364A),.A2(g4679A),.A1(g1215A));
AND2_X1 U_g9649A (.ZN(g9649A),.A2(g9205A),.A1(g916A));
AND2_X1 U_g5795A (.ZN(g5795A),.A2(g5261A),.A1(g1543A));
AND2_X1 U_g5737A (.ZN(g5737A),.A2(FE_OFN321_g5261A),.A1(g1524A));
AND2_X1 U_g6841A (.ZN(g6841A),.A2(FE_OFN180_g5354A),.A1(g1400A));
AND2_X1 U_g4054A (.ZN(g4054A),.A2(g2774A),.A1(g1753A));
AND2_X1 U_g6345A (.ZN(g6345A),.A2(FE_OFN346_g4381A),.A1(g5823A));
AND2_X1 U_g11391A (.ZN(g11391A),.A2(g7914A),.A1(g11275A));
AND2_X1 U_g9851A (.ZN(g9851A),.A2(g9764A),.A1(g296A));
AND2_X1 U_g6763A (.ZN(g6763A),.A2(g4381A),.A1(g5802A));
AND2_X1 U_g4770A (.ZN(g4770A),.A2(FE_OFN300_g4002A),.A1(g416A));
AND3_X1 U_I16142A (.ZN(I16142A),.A3(g10507A),.A2(g10509A),.A1(g10511A));
AND2_X1 U_g9698A (.ZN(g9698A),.A2(FE_OFN63_g9474A),.A1(g1571A));
AND2_X1 U_g4725A (.ZN(g4725A),.A2(FE_OFN347_g3914A),.A1(g1032A));
AND2_X1 U_g5477A (.ZN(g5477A),.A2(FE_OFN333_g4294A),.A1(g1887A));
AND2_X1 U_g9964A (.ZN(g9964A),.A2(g9536A),.A1(g9954A));
AND2_X1 U_g5523A (.ZN(g5523A),.A2(g4290A),.A1(g1663A));
AND2_X1 U_g4553A (.ZN(g4553A),.A2(g4002A),.A1(g435A));
AND2_X1 U_g8550A (.ZN(g8550A),.A2(FE_OFN330_g7638A),.A1(g8402A));
AND2_X1 U_g8845A (.ZN(g8845A),.A2(FE_OFN328_g8709A),.A1(g8611A));
AND2_X1 U_g2081A (.ZN(g2081A),.A2(g928A),.A1(g932A));
AND2_X1 U_g6359A (.ZN(g6359A),.A2(FE_OFN320_g5361A),.A1(g281A));
AND2_X1 U_g11586A (.ZN(g11586A),.A2(g11539A),.A1(g1324A));
AND2_X1 U_g11007A (.ZN(g11007A),.A2(FE_OFN13_g10702A),.A1(g5147A));
AND2_X1 U_g5104A (.ZN(g5104A),.A2(g4608A),.A1(g1796A));
AND2_X1 U_g5099A (.ZN(g5099A),.A2(FE_OFN141_g3829A),.A1(g4821A));
AND2_X1 U_g6757A (.ZN(g6757A),.A2(g5919A),.A1(g143A));
AND2_X1 U_g5499A (.ZN(g5499A),.A2(g4679A),.A1(g1627A));
AND2_X1 U_g4389A (.ZN(g4389A),.A2(g3092A),.A1(g3529A));
AND2_X1 U_g6416A (.ZN(g6416A),.A2(FE_OFN217_g5013A),.A1(g3497A));
AND2_X1 U_g9720A (.ZN(g9720A),.A2(g9490A),.A1(g1546A));
AND2_X1 U_g4990A (.ZN(g4990A),.A2(FE_OFN147_g4682A),.A1(g1444A));
AND2_X1 U_g9619A (.ZN(g9619A),.A2(g9010A),.A1(g940A));
AND4_X1 U_I6630A (.ZN(I6630A),.A4(FE_OFN253_g1786A),.A3(FE_OFN236_g1776A),.A2(FE_OFN247_g1771A),.A1(g2677A));
AND2_X1 U_g6047A (.ZN(g6047A),.A2(g4977A),.A1(g2017A));
AND2_X1 U_g9652A (.ZN(g9652A),.A2(FE_OFN39_g9223A),.A1(g953A));
AND3_X1 U_g10515A (.ZN(g10515A),.A3(I16142A),.A2(g10469A),.A1(g10505A));
AND2_X1 U_g9843A (.ZN(g9843A),.A2(g9519A),.A1(g9711A));
AND2_X1 U_g5273A (.ZN(g5273A),.A2(g4776A),.A1(g1074A));
AND2_X1 U_g11465A (.ZN(g11465A),.A2(FE_OFN100_g4421A),.A1(g11232A));
AND2_X1 U_g5044A (.ZN(g5044A),.A2(g1918A),.A1(g4348A));
AND2_X1 U_g11237A (.ZN(g11237A),.A2(g11111A),.A1(g4548A));
AND2_X1 U_g9834A (.ZN(g9834A),.A2(FE_OFN34_g9785A),.A1(g9731A));
AND2_X1 U_g6654A (.ZN(g6654A),.A2(FE_OFN282_g6165A),.A1(g363A));
AND2_X1 U_g5444A (.ZN(g5444A),.A2(FE_OFN290_g4880A),.A1(g1041A));
AND2_X1 U_g3714A (.ZN(g3714A),.A2(g2299A),.A1(g1690A));
AND2_X1 U_g11340A (.ZN(g11340A),.A2(g4285A),.A1(g11285A));
AND2_X1 U_g9598A (.ZN(g9598A),.A2(g9274A),.A1(g119A));
AND2_X1 U_g8097A (.ZN(g8097A),.A2(g7852A),.A1(g5477A));
AND2_X1 U_g8726A (.ZN(g8726A),.A2(g7913A),.A1(g8221A));
AND2_X1 U_g6880A (.ZN(g6880A),.A2(g6557A),.A1(g4816A));
AND2_X1 U_g4338A (.ZN(g4338A),.A2(FE_OFN351_g3913A),.A1(g1157A));
AND2_X1 U_g5543A (.ZN(g5543A),.A2(FE_OFN322_g4449A),.A1(g2979A));
AND3_X1 U_g8960A (.ZN(g8960A),.A3(g8828A),.A2(FE_OFN95_g2216A),.A1(g8085A));
AND2_X1 U_g4109A (.ZN(g4109A),.A2(g3287A),.A1(g806A));
AND2_X1 U_g10759A (.ZN(g10759A),.A2(g10556A),.A1(g10557A));
AND2_X1 U_g9938A (.ZN(g9938A),.A2(FE_OFN67_g9367A),.A1(g9917A));
AND2_X1 U_g10758A (.ZN(g10758A),.A2(FE_OFN293_g3015A),.A1(g10652A));
AND2_X1 U_g4759A (.ZN(g4759A),.A2(FE_OFN300_g4002A),.A1(g406A));
AND2_X1 U_g9909A (.ZN(g9909A),.A2(FE_OFN33_g9454A),.A1(g9891A));
AND2_X1 U_g7127A (.ZN(g7127A),.A2(g2241A),.A1(g6663A));
AND2_X1 U_g11165A (.ZN(g11165A),.A2(FE_OFN13_g10702A),.A1(g476A));
AND2_X1 U_g6234A (.ZN(g6234A),.A2(FE_OFN306_g5128A),.A1(g1424A));
AND2_X1 U_g6328A (.ZN(g6328A),.A2(FE_OFN115_g4807A),.A1(g1260A));
AND2_X1 U_g8401A (.ZN(g8401A),.A2(g8146A),.A1(g677A));
AND2_X1 U_g11006A (.ZN(g11006A),.A2(FE_OFN18_g10702A),.A1(g5125A));
AND2_X1 U_g4865A (.ZN(g4865A),.A2(FE_OFN297_g3015A),.A1(g1080A));
AND2_X1 U_g4715A (.ZN(g4715A),.A2(FE_OFN297_g3015A),.A1(g1077A));
AND3_X1 U_g4604A (.ZN(g4604A),.A3(g2325A),.A2(g3753A),.A1(g3056A));
AND2_X1 U_g5513A (.ZN(g5513A),.A2(g3906A),.A1(g1675A));
AND2_X1 U_g11222A (.ZN(g11222A),.A2(FE_OFN279_g11157A),.A1(g965A));
AND2_X1 U_g4498A (.ZN(g4498A),.A2(FE_OFN302_g3913A),.A1(g1145A));
AND2_X1 U_g6554A (.ZN(g6554A),.A2(g5808A),.A1(g96A));
AND2_X1 U_g7732A (.ZN(g7732A),.A2(FE_OFN226_g3880A),.A1(g5803A));
AND2_X1 U_g9586A (.ZN(g9586A),.A2(FE_OFN53_g9173A),.A1(g1346A));
AND3_X1 U_g5178A (.ZN(g5178A),.A3(g4104A),.A2(FE_OFN223_g4401A),.A1(g2047A));
AND2_X1 U_g4584A (.ZN(g4584A),.A2(g1857A),.A1(g3710A));
AND2_X1 U_g7472A (.ZN(g7472A),.A2(g61A),.A1(FE_OFN83_g2176A));
AND2_X1 U_g11253A (.ZN(g11253A),.A2(g11083A),.A1(g981A));
AND2_X1 U_g5182A (.ZN(g5182A),.A2(FE_OFN303_g4678A),.A1(g1240A));
AND2_X1 U_g9860A (.ZN(g9860A),.A2(g9778A),.A1(g1598A));
AND2_X1 U_g11600A (.ZN(g11600A),.A2(g11575A),.A1(g1346A));
AND2_X1 U_g9710A (.ZN(g9710A),.A2(FE_OFN63_g9474A),.A1(g1586A));
AND2_X1 U_g9645A (.ZN(g9645A),.A2(FE_OFN51_g9111A),.A1(g1203A));
AND2_X1 U_g11236A (.ZN(g11236A),.A2(g11111A),.A1(g4537A));
AND2_X1 U_g4162A (.ZN(g4162A),.A2(g1845A),.A1(g3106A));
AND2_X1 U_g6090A (.ZN(g6090A),.A2(g5627A),.A1(g553A));
AND2_X1 U_g9691A (.ZN(g9691A),.A2(g9432A),.A1(g269A));
AND2_X1 U_g11372A (.ZN(g11372A),.A2(g4285A),.A1(g11316A));
AND2_X1 U_g6823A (.ZN(g6823A),.A2(g5354A),.A1(g1368A));
AND2_X1 U_g11175A (.ZN(g11175A),.A2(FE_OFN20_g10702A),.A1(g501A));
AND2_X1 U_g8068A (.ZN(g8068A),.A2(FE_OFN198_g7697A),.A1(g664A));
AND2_X1 U_g9607A (.ZN(g9607A),.A2(g9274A),.A1(g12A));
AND2_X1 U_g9962A (.ZN(g9962A),.A2(FE_OFN280_g9536A),.A1(g9952A));
AND2_X1 U_g6348A (.ZN(g6348A),.A2(FE_OFN320_g5361A),.A1(g296A));
AND2_X1 U_g9659A (.ZN(g9659A),.A2(FE_OFN39_g9223A),.A1(g956A));
AND2_X1 U_g9358A (.ZN(g9358A),.A2(FE_OFN47_g9151A),.A1(g1318A));
AND2_X1 U_g3104A (.ZN(g3104A),.A2(I6317A),.A1(I6316A));
AND2_X1 U_g4486A (.ZN(g4486A),.A2(g4679A),.A1(g1711A));
AND2_X1 U_g9587A (.ZN(g9587A),.A2(g8995A),.A1(g892A));
AND2_X1 U_g5632A (.ZN(g5632A),.A2(I5435A),.A1(g1636A));
AND2_X4 U_g9111A (.ZN(g9111A),.A2(FE_OFN276_g48A),.A1(g8965A));
AND2_X1 U_g4881A (.ZN(g4881A),.A2(FE_OFN347_g3914A),.A1(g991A));
AND2_X1 U_g11209A (.ZN(g11209A),.A2(FE_OFN79_g8700A),.A1(g10712A));
AND2_X1 U_g8848A (.ZN(g8848A),.A2(FE_OFN328_g8709A),.A1(g8715A));
AND2_X1 U_g4070A (.ZN(g4070A),.A2(g2330A),.A1(g3263A));
AND2_X1 U_g6463A (.ZN(g6463A),.A2(I9237A),.A1(FE_OFN277_g48A));
AND4_X1 U_I5689A (.ZN(I5689A),.A4(g1432A),.A3(g1428A),.A2(g1424A),.A1(g1419A));
AND2_X1 U_g7820A (.ZN(g7820A),.A2(FE_OFN209_g6863A),.A1(g1896A));
AND2_X1 U_g11021A (.ZN(g11021A),.A2(FE_OFN7_g10702A),.A1(g448A));
AND2_X1 U_g5917A (.ZN(g5917A),.A2(g85A),.A1(g1044A));
AND2_X1 U_g6619A (.ZN(g6619A),.A2(FE_OFN97_I8869A),.A1(g49A));
AND2_X1 U_g6318A (.ZN(g6318A),.A2(FE_OFN118_g4807A),.A1(g1300A));
AND2_X1 U_g6872A (.ZN(g6872A),.A2(FE_OFN213_g6003A),.A1(g1896A));
AND2_X1 U_g11320A (.ZN(g11320A),.A2(g4379A),.A1(g11201A));
AND2_X1 U_g10514A (.ZN(g10514A),.A2(FE_OFN370_g4525A),.A1(g10489A));
AND2_X1 U_g4006A (.ZN(g4006A),.A2(FE_OFN266_g18A),.A1(g201A));
AND2_X1 U_g9853A (.ZN(g9853A),.A2(g9764A),.A1(g299A));
AND2_X1 U_g11274A (.ZN(g11274A),.A2(g11199A),.A1(g4771A));
AND2_X1 U_g6193A (.ZN(g6193A),.A2(FE_OFN306_g5128A),.A1(g1419A));
AND2_X1 U_g8119A (.ZN(g8119A),.A2(FE_OFN207_g6863A),.A1(g5526A));
AND2_X1 U_g9420A (.ZN(g9420A),.A2(FE_OFN50_g9030A),.A1(g1747A));
AND2_X1 U_g5233A (.ZN(g5233A),.A2(g4492A),.A1(FE_OFN252_g1791A));
AND2_X1 U_g7581A (.ZN(g7581A),.A2(g5420A),.A1(g7092A));
AND2_X1 U_g6549A (.ZN(g6549A),.A2(g5808A),.A1(g95A));
AND2_X1 U_g11464A (.ZN(g11464A),.A2(FE_OFN100_g4421A),.A1(g11231A));
AND2_X1 U_g4801A (.ZN(g4801A),.A2(FE_OFN307_g4010A),.A1(g516A));
AND2_X1 U_g6834A (.ZN(g6834A),.A2(FE_OFN178_g5354A),.A1(g1365A));
AND2_X1 U_g4487A (.ZN(g4487A),.A2(g3906A),.A1(g1718A));
AND2_X1 U_g2939A (.ZN(g2939A),.A2(g1687A),.A1(FE_OFN241_g1690A));
AND2_X1 U_g7060A (.ZN(g7060A),.A2(g5521A),.A1(g6739A));
AND2_X1 U_g5770A (.ZN(g5770A),.A2(g5128A),.A1(g3585A));
AND2_X1 U_g5725A (.ZN(g5725A),.A2(FE_OFN353_g5117A),.A1(g1580A));
AND2_X1 U_g11641A (.ZN(g11641A),.A2(g7897A),.A1(g11615A));
AND2_X1 U_g2544A (.ZN(g2544A),.A2(g1336A),.A1(g1341A));
AND2_X1 U_g11292A (.ZN(g11292A),.A2(g4379A),.A1(g11252A));
AND2_X1 U_g5532A (.ZN(g5532A),.A2(g4273A),.A1(g1681A));
AND2_X1 U_g11153A (.ZN(g11153A),.A2(g10788A),.A1(g3771A));
AND2_X1 U_g9905A (.ZN(g9905A),.A2(g9680A),.A1(g9872A));
AND2_X1 U_g7739A (.ZN(g7739A),.A2(g3880A),.A1(g5820A));
AND2_X1 U_g6321A (.ZN(g6321A),.A2(FE_OFN118_g4807A),.A1(g1284A));
AND2_X1 U_g8386A (.ZN(g8386A),.A2(g8220A),.A1(g5257A));
AND3_X1 U_g8975A (.ZN(g8975A),.A3(FE_OFN73_g8858A),.A2(FE_OFN281_g2216A),.A1(g8089A));
AND2_X1 U_g2306A (.ZN(g2306A),.A2(g1218A),.A1(g1223A));
AND2_X1 U_g6625A (.ZN(g6625A),.A2(g6081A),.A1(g1218A));
AND2_X1 U_g7937A (.ZN(g7937A),.A2(FE_OFN292_g3015A),.A1(g5274A));
AND2_X2 U_g10788A (.ZN(g10788A),.A2(g10702A),.A1(g8303A));
AND2_X1 U_g10325A (.ZN(g10325A),.A2(FE_OFN352_g109A),.A1(I15503A));
AND2_X1 U_g8170A (.ZN(g8170A),.A2(FE_OFN89_I11360A),.A1(g36A));
AND2_X1 U_g5706A (.ZN(g5706A),.A2(FE_OFN315_g5117A),.A1(g1574A));
AND2_X1 U_g2756A (.ZN(g2756A),.A2(g2081A),.A1(g936A));
AND2_X1 U_g8821A (.ZN(g8821A),.A2(FE_OFN328_g8709A),.A1(g8643A));
AND2_X1 U_g10946A (.ZN(g10946A),.A2(FE_OFN9_g10702A),.A1(g5225A));
AND2_X1 U_g4169A (.ZN(g4169A),.A2(g3060A),.A1(FE_OFN237_g1806A));
AND2_X1 U_g5029A (.ZN(g5029A),.A2(FE_OFN288_g4263A),.A1(g1077A));
AND2_X1 U_g11164A (.ZN(g11164A),.A2(FE_OFN13_g10702A),.A1(g3513A));
AND2_X1 U_g4007A (.ZN(g4007A),.A2(g2276A),.A1(FE_OFN247_g1771A));
AND2_X1 U_g4059A (.ZN(g4059A),.A2(g2774A),.A1(g1756A));
AND2_X1 U_g4868A (.ZN(g4868A),.A2(FE_OFN347_g3914A),.A1(g1027A));
AND2_X1 U_g5675A (.ZN(g5675A),.A2(FE_OFN365_g5361A),.A1(g131A));
AND2_X1 U_g4718A (.ZN(g4718A),.A2(g3943A),.A1(g650A));
AND2_X1 U_g10682A (.ZN(g10682A),.A2(FE_OFN136_g3863A),.A1(g10381A));
AND2_X1 U_g6687A (.ZN(g6687A),.A2(I9326A),.A1(g92A));
AND2_X1 U_g7704A (.ZN(g7704A),.A2(FE_OFN191_g6488A),.A1(g682A));
AND2_X1 U_g4582A (.ZN(g4582A),.A2(g4010A),.A1(g525A));
AND2_X1 U_g4261A (.ZN(g4261A),.A2(FE_OFN347_g3914A),.A1(g1019A));
AND2_X1 U_g3422A (.ZN(g3422A),.A2(FE_OFN324_g18A),.A1(g225A));
AND2_X1 U_g5745A (.ZN(g5745A),.A2(FE_OFN321_g5261A),.A1(g1549A));
AND2_X1 U_g8387A (.ZN(g8387A),.A2(g8220A),.A1(g5258A));
AND2_X1 U_g7954A (.ZN(g7954A),.A2(g7512A),.A1(g49A));
AND2_X1 U_g11283A (.ZN(g11283A),.A2(g11239A),.A1(g4804A));
AND2_X1 U_g8461A (.ZN(g8461A),.A2(FE_OFN210_g7246A),.A1(g8298A));
AND2_X1 U_g10760A (.ZN(g10760A),.A2(g10554A),.A1(g10555A));
AND2_X1 U_g11492A (.ZN(g11492A),.A2(g4807A),.A1(g11480A));
AND3_X1 U_g7032A (.ZN(g7032A),.A3(I7048A),.A2(g6626A),.A1(g109A));
AND2_X4 U_g9151A (.ZN(g9151A),.A2(FE_OFN276_g48A),.A1(g8967A));
AND2_X1 U_g6341A (.ZN(g6341A),.A2(FE_OFN319_g5361A),.A1(g272A));
AND2_X1 U_g10506A (.ZN(g10506A),.A2(FE_OFN241_g1690A),.A1(g10007A));
AND2_X1 U_g9648A (.ZN(g9648A),.A2(FE_OFN62_g9274A),.A1(g16A));
AND2_X1 U_g7453A (.ZN(g7453A),.A2(g52A),.A1(FE_OFN86_g2176A));
AND2_X1 U_g6525A (.ZN(g6525A),.A2(FE_OFN343_I5565A),.A1(g5995A));
AND2_X1 U_g6645A (.ZN(g6645A),.A2(FE_OFN97_I8869A),.A1(g67A));
AND2_X1 U_g5707A (.ZN(g5707A),.A2(FE_OFN353_g5117A),.A1(g1595A));
AND2_X1 U_g8046A (.ZN(g8046A),.A2(FE_OFN305_g5151A),.A1(g7548A));
AND2_X1 U_g11091A (.ZN(g11091A),.A2(FE_OFN4_g10950A),.A1(g833A));
AND2_X1 U_g11174A (.ZN(g11174A),.A2(FE_OFN21_g10702A),.A1(g496A));
AND2_X4 U_g9010A (.ZN(g9010A),.A2(g8930A),.A1(FE_OFN277_g48A));
AND2_X1 U_g8403A (.ZN(g8403A),.A2(g8220A),.A1(g5276A));
AND2_X1 U_g5201A (.ZN(g5201A),.A2(g4678A),.A1(g1250A));
AND2_X1 U_g8841A (.ZN(g8841A),.A2(FE_OFN328_g8709A),.A1(g8605A));
AND2_X1 U_g6879A (.ZN(g6879A),.A2(FE_OFN213_g6003A),.A1(g1914A));
AND2_X2 U_g8763A (.ZN(g8763A),.A2(g8451A),.A1(I9880A));
AND2_X1 U_g4502A (.ZN(g4502A),.A2(g3938A),.A1(g2031A));
AND2_X1 U_g9839A (.ZN(g9839A),.A2(g9747A),.A1(g9702A));
AND2_X1 U_g6358A (.ZN(g6358A),.A2(FE_OFN346_g4381A),.A1(g5841A));
AND2_X1 U_g5575A (.ZN(g5575A),.A2(FE_OFN367_g3521A),.A1(g1618A));
AND2_X1 U_g4940A (.ZN(g4940A),.A2(FE_OFN310_g4336A),.A1(g1984A));
AND2_X1 U_g8107A (.ZN(g8107A),.A2(g7852A),.A1(g5502A));
AND2_X1 U_g10240A (.ZN(g10240A),.A2(g9082A),.A1(g9974A));
AND2_X1 U_g11192A (.ZN(g11192A),.A2(g10927A),.A1(g4759A));
AND2_X1 U_g9618A (.ZN(g9618A),.A2(g9205A),.A1(g910A));
AND2_X1 U_g5539A (.ZN(g5539A),.A2(g4273A),.A1(g1684A));
AND2_X1 U_g8416A (.ZN(g8416A),.A2(FE_OFN187_g7638A),.A1(g731A));
AND2_X1 U_g9693A (.ZN(g9693A),.A2(FE_OFN59_g9432A),.A1(g275A));
AND2_X1 U_g11553A (.ZN(g11553A),.A2(g11519A),.A1(g1771A));
AND2_X1 U_g8047A (.ZN(g8047A),.A2(FE_OFN177_g5919A),.A1(g7557A));
AND2_X1 U_g5268A (.ZN(g5268A),.A2(g4263A),.A1(g1098A));
AND2_X1 U_g9555A (.ZN(g9555A),.A2(FE_OFN325_g18A),.A1(g9107A));
AND2_X1 U_g6180A (.ZN(g6180A),.A2(g5128A),.A1(g1453A));
AND2_X1 U_g6832A (.ZN(g6832A),.A2(FE_OFN179_g5354A),.A1(g1383A));
AND2_X1 U_g10633A (.ZN(g10633A),.A2(g3829A),.A1(g10381A));
AND2_X1 U_g7894A (.ZN(g7894A),.A2(FE_OFN366_g3521A),.A1(g5317A));
AND2_X1 U_g8654A (.ZN(g8654A),.A2(FE_OFN348_g3015A),.A1(g8266A));
AND2_X1 U_g9621A (.ZN(g9621A),.A2(FE_OFN46_g9125A),.A1(g1179A));
AND2_X1 U_g6794A (.ZN(g6794A),.A2(FE_OFN346_g4381A),.A1(g5819A));
AND2_X1 U_g9313A (.ZN(g9313A),.A2(FE_OFN275_g48A),.A1(g8876A));
AND2_X1 U_g3412A (.ZN(g3412A),.A2(g18A),.A1(g219A));
AND2_X1 U_g7661A (.ZN(g7661A),.A2(g2251A),.A1(g7127A));
AND3_X1 U_g2800A (.ZN(g2800A),.A3(g591A),.A2(g2369A),.A1(g2399A));
AND2_X1 U_g3706A (.ZN(g3706A),.A2(g3268A),.A1(g471A));
AND2_X1 U_g9908A (.ZN(g9908A),.A2(FE_OFN33_g9454A),.A1(g9760A));
AND2_X1 U_g3429A (.ZN(g3429A),.A2(g18A),.A1(g231A));
AND2_X1 U_g6628A (.ZN(g6628A),.A2(FE_OFN282_g6165A),.A1(g351A));
AND2_X1 U_g5470A (.ZN(g5470A),.A2(g4880A),.A1(g1044A));
AND2_X1 U_g7526A (.ZN(g7526A),.A2(g73A),.A1(FE_OFN87_g2176A));
AND2_X1 U_g5897A (.ZN(g5897A),.A2(g5354A),.A1(g2204A));
AND2_X1 U_g5025A (.ZN(g5025A),.A2(FE_OFN153_g4640A),.A1(g1482A));
AND2_X1 U_g6204A (.ZN(g6204A),.A2(FE_OFN200_g4921A),.A1(g3738A));
AND2_X1 U_g4048A (.ZN(g4048A),.A2(g2774A),.A1(g1750A));
AND3_X1 U_g8935A (.ZN(g8935A),.A3(g8849A),.A2(FE_OFN95_g2216A),.A1(g8106A));
AND2_X1 U_g3281A (.ZN(g3281A),.A2(g2525A),.A1(g766A));
AND2_X1 U_g9593A (.ZN(g9593A),.A2(FE_OFN42_g9205A),.A1(g898A));
AND2_X1 U_g4827A (.ZN(g4827A),.A2(FE_OFN324_g18A),.A1(g213A));
AND2_X1 U_g10701A (.ZN(g10701A),.A2(g10500A),.A1(g10501A));
AND2_X1 U_g10777A (.ZN(g10777A),.A2(g3015A),.A1(g10733A));
AND2_X1 U_g8130A (.ZN(g8130A),.A2(g7952A),.A1(g1936A));
AND2_X1 U_g9965A (.ZN(g9965A),.A2(FE_OFN280_g9536A),.A1(g9955A));
AND2_X1 U_g3684A (.ZN(g3684A),.A2(g3015A),.A1(g1710A));
AND2_X1 U_g11213A (.ZN(g11213A),.A2(FE_OFN279_g11157A),.A1(g947A));
AND2_X1 U_g5006A (.ZN(g5006A),.A2(FE_OFN154_g4640A),.A1(g1462A));
AND2_X1 U_g9933A (.ZN(g9933A),.A2(g9624A),.A1(g9912A));
AND2_X1 U_g8554A (.ZN(g8554A),.A2(FE_OFN330_g7638A),.A1(g8407A));
AND2_X1 U_g9641A (.ZN(g9641A),.A2(g9205A),.A1(g913A));
AND2_X1 U_g6123A (.ZN(g6123A),.A2(FE_OFN310_g4336A),.A1(g3662A));
AND2_X1 U_g6323A (.ZN(g6323A),.A2(FE_OFN116_g4807A),.A1(g1235A));
AND2_X1 U_g10766A (.ZN(g10766A),.A2(FE_OFN131_g3015A),.A1(g10646A));
AND2_X1 U_g6666A (.ZN(g6666A),.A2(g5836A),.A1(g89A));
AND2_X1 U_g4994A (.ZN(g4994A),.A2(FE_OFN154_g4640A),.A1(g1504A));
AND2_X1 U_g5755A (.ZN(g5755A),.A2(FE_OFN179_g5354A),.A1(g5103A));
AND2_X1 U_g11592A (.ZN(g11592A),.A2(g11561A),.A1(g3717A));
AND2_X1 U_g6351A (.ZN(g6351A),.A2(g48A),.A1(I9237A));
AND2_X1 U_g6875A (.ZN(g6875A),.A2(FE_OFN213_g6003A),.A1(g1905A));
AND2_X1 U_g4816A (.ZN(g4816A),.A2(g2336A),.A1(g4070A));
AND2_X1 U_g9658A (.ZN(g9658A),.A2(g9240A),.A1(g947A));
AND2_X1 U_g6530A (.ZN(g6530A),.A2(FE_OFN141_g3829A),.A1(g6207A));
AND2_X1 U_g8366A (.ZN(g8366A),.A2(g7265A),.A1(g8199A));
AND2_X1 U_g9835A (.ZN(g9835A),.A2(FE_OFN34_g9785A),.A1(g9735A));
AND2_X1 U_g6655A (.ZN(g6655A),.A2(I9326A),.A1(g88A));
AND3_X1 U_g5445A (.ZN(g5445A),.A3(g109A),.A2(g3875A),.A1(FE_OFN184_I7048A));
AND2_X1 U_g5173A (.ZN(g5173A),.A2(g4671A),.A1(g1110A));
AND2_X1 U_g7970A (.ZN(g7970A),.A2(g7438A),.A1(g7384A));
AND2_X1 U_g3098A (.ZN(g3098A),.A2(g2198A),.A1(g2331A));
AND2_X1 U_g5491A (.ZN(g5491A),.A2(g4289A),.A1(g1624A));
AND2_X1 U_g9271A (.ZN(g9271A),.A2(g8949A),.A1(g6109A));
AND2_X1 U_g11152A (.ZN(g11152A),.A2(g10883A),.A1(g369A));
AND2_X1 U_g9611A (.ZN(g9611A),.A2(g9010A),.A1(g936A));
AND2_X1 U_g6410A (.ZN(g6410A),.A2(FE_OFN217_g5013A),.A1(g2804A));
AND2_X1 U_g10451A (.ZN(g10451A),.A2(g2024A),.A1(g10444A));
AND2_X1 U_g4397A (.ZN(g4397A),.A2(g639A),.A1(g3475A));
AND2_X1 U_g7224A (.ZN(g7224A),.A2(g6447A),.A1(g5398A));
AND2_X1 U_g5602A (.ZN(g5602A),.A2(FE_OFN357_g3521A),.A1(g1624A));
AND2_X2 U_g4421A (.ZN(g4421A),.A2(g750A),.A1(g2057A));
AND2_X1 U_g6884A (.ZN(g6884A),.A2(g6557A),.A1(g5569A));
AND2_X1 U_g6839A (.ZN(g6839A),.A2(FE_OFN180_g5354A),.A1(g1397A));
AND3_X1 U_g8964A (.ZN(g8964A),.A3(g8849A),.A2(FE_OFN92_g2216A),.A1(g8255A));
AND2_X1 U_g8260A (.ZN(g8260A),.A2(g7907A),.A1(g940A));
AND2_X1 U_g11413A (.ZN(g11413A),.A2(g10679A),.A1(g11217A));
AND2_X1 U_g4950A (.ZN(g4950A),.A2(FE_OFN146_g4682A),.A1(g1415A));
AND2_X1 U_g5535A (.ZN(g5535A),.A2(FE_OFN366_g3521A),.A1(g572A));
AND2_X1 U_g7277A (.ZN(g7277A),.A2(g731A),.A1(g6772A));
AND2_X1 U_g8463A (.ZN(g8463A),.A2(FE_OFN211_g7246A),.A1(g8301A));
AND2_X1 U_g3268A (.ZN(g3268A),.A2(g2511A),.A1(FE_OFN248_g466A));
AND2_X1 U_g10785A (.ZN(g10785A),.A2(g4467A),.A1(g10728A));
AND2_X1 U_g6618A (.ZN(g6618A),.A2(FE_OFN219_g5557A),.A1(g658A));
AND2_X1 U_g6235A (.ZN(g6235A),.A2(g5613A),.A1(g569A));
AND2_X1 U_g10950A (.ZN(g10950A),.A2(g6355A),.A1(g10788A));
AND2_X1 U_g4723A (.ZN(g4723A),.A2(g627A),.A1(g3626A));
AND2_X1 U_g8720A (.ZN(g8720A),.A2(g7905A),.A1(g8206A));
AND2_X1 U_g6693A (.ZN(g6693A),.A2(I9326A),.A1(g93A));
AND2_X1 U_g11020A (.ZN(g11020A),.A2(FE_OFN7_g10702A),.A1(g452A));
AND2_X1 U_g11583A (.ZN(g11583A),.A2(g11539A),.A1(g1314A));
AND2_X1 U_g8118A (.ZN(g8118A),.A2(g7949A),.A1(g1900A));
AND2_X1 U_g8167A (.ZN(g8167A),.A2(FE_OFN89_I11360A),.A1(g33A));
AND2_X1 U_g6334A (.ZN(g6334A),.A2(FE_OFN180_g5354A),.A1(g1389A));
AND2_X1 U_g7892A (.ZN(g7892A),.A2(g3814A),.A1(g5308A));
AND2_X1 U_g8652A (.ZN(g8652A),.A2(FE_OFN119_g3015A),.A1(g8264A));
AND2_X1 U_g5721A (.ZN(g5721A),.A2(FE_OFN353_g5117A),.A1(g1577A));
AND2_X1 U_g10367A (.ZN(g10367A),.A2(FE_OFN234_g2024A),.A1(g10362A));
AND2_X1 U_g9901A (.ZN(g9901A),.A2(FE_OFN69_g9392A),.A1(g9719A));
AND2_X1 U_g6792A (.ZN(g6792A),.A2(FE_OFN319_g5361A),.A1(g290A));
AND2_X1 U_g11282A (.ZN(g11282A),.A2(g11203A),.A1(g4801A));
AND2_X1 U_g7945A (.ZN(g7945A),.A2(g7473A),.A1(g67A));
AND3_X1 U_g8971A (.ZN(g8971A),.A3(FE_OFN73_g8858A),.A2(FE_OFN281_g2216A),.A1(g8081A));
AND2_X1 U_g11302A (.ZN(g11302A),.A2(g11243A),.A1(g4582A));
AND2_X1 U_g4585A (.ZN(g4585A),.A2(g4010A),.A1(g521A));
AND2_X1 U_g6621A (.ZN(g6621A),.A2(I8869A),.A1(g52A));
AND2_X1 U_g5502A (.ZN(g5502A),.A2(FE_OFN333_g4294A),.A1(g1932A));
AND2_X1 U_g11105A (.ZN(g11105A),.A2(g10937A),.A1(g3634A));
AND2_X1 U_g7709A (.ZN(g7709A),.A2(FE_OFN322_g4449A),.A1(g5942A));
AND2_X1 U_g8598A (.ZN(g8598A),.A2(FE_OFN210_g7246A),.A1(g8471A));
AND2_X1 U_g7140A (.ZN(g7140A),.A2(g6716A),.A1(g5221A));
AND2_X1 U_g9600A (.ZN(g9600A),.A2(FE_OFN42_g9205A),.A1(g904A));
AND2_X1 U_g9864A (.ZN(g9864A),.A2(g9778A),.A1(g1604A));
AND2_X1 U_g11640A (.ZN(g11640A),.A2(g7897A),.A1(g11613A));
AND2_X1 U_g5188A (.ZN(g5188A),.A2(g794A),.A1(g798A));
AND2_X1 U_g7435A (.ZN(g7435A),.A2(g6403A),.A1(g7260A));
AND2_X1 U_g7876A (.ZN(g7876A),.A2(FE_OFN366_g3521A),.A1(g5278A));
AND2_X1 U_g5030A (.ZN(g5030A),.A2(FE_OFN303_g4678A),.A1(g1280A));
AND2_X1 U_g4058A (.ZN(g4058A),.A2(FE_OFN224_g2276A),.A1(FE_OFN252_g1791A));
AND2_X1 U_g6776A (.ZN(g6776A),.A2(FE_OFN111_g3914A),.A1(g5809A));
AND2_X1 U_g4890A (.ZN(g4890A),.A2(g4739A),.A1(g630A));
AND2_X1 U_g2525A (.ZN(g2525A),.A2(g758A),.A1(g762A));
AND2_X1 U_g10301A (.ZN(g10301A),.A2(g10025A),.A1(g8700A));
AND2_X1 U_g4505A (.ZN(g4505A),.A2(FE_OFN287_g3586A),.A1(g354A));
AND2_X1 U_g9623A (.ZN(g9623A),.A2(FE_OFN62_g9274A),.A1(g17A));
AND2_X1 U_g10739A (.ZN(g10739A),.A2(g3368A),.A1(g10676A));
AND2_X1 U_g11027A (.ZN(g11027A),.A2(FE_OFN17_g10702A),.A1(g391A));
AND2_X1 U_g10738A (.ZN(g10738A),.A2(FE_OFN131_g3015A),.A1(g10599A));
AND2_X1 U_g8687A (.ZN(g8687A),.A2(FE_OFN189_g7638A),.A1(g8558A));
AND2_X1 U_g6360A (.ZN(g6360A),.A2(FE_OFN319_g5361A),.A1(g302A));
AND2_X1 U_g9871A (.ZN(g9871A),.A2(g9802A),.A1(g1564A));
AND2_X1 U_g5108A (.ZN(g5108A),.A2(g4608A),.A1(g1801A));
AND2_X1 U_g11248A (.ZN(g11248A),.A2(g11083A),.A1(g976A));
AND2_X1 U_g4992A (.ZN(g4992A),.A2(FE_OFN147_g4682A),.A1(g1407A));
AND2_X1 U_g11552A (.ZN(g11552A),.A2(FE_OFN27_g11519A),.A1(g2677A));
AND2_X1 U_g9651A (.ZN(g9651A),.A2(g9240A),.A1(g944A));
AND2_X1 U_g11204A (.ZN(g11204A),.A2(g11083A),.A1(g971A));
AND2_X1 U_g7824A (.ZN(g7824A),.A2(FE_OFN206_g6863A),.A1(g1932A));
AND2_X1 U_g4480A (.ZN(g4480A),.A2(FE_OFN302_g3913A),.A1(g1133A));
AND2_X1 U_g6179A (.ZN(g6179A),.A2(g5354A),.A1(g5115A));
AND2_X1 U_g7590A (.ZN(g7590A),.A2(g5420A),.A1(g7102A));
AND2_X1 U_g9384A (.ZN(g9384A),.A2(g9223A),.A1(g968A));
AND2_X1 U_g3407A (.ZN(g3407A),.A2(FE_OFN352_g109A),.A1(g2561A));
AND2_X1 U_g9838A (.ZN(g9838A),.A2(g9754A),.A1(g9700A));
AND2_X1 U_g10661A (.ZN(g10661A),.A2(FE_OFN119_g3015A),.A1(g10594A));
AND2_X1 U_g11380A (.ZN(g11380A),.A2(g4285A),.A1(g11321A));
AND3_X1 U_g8879A (.ZN(g8879A),.A3(FE_OFN73_g8858A),.A2(FE_OFN281_g2216A),.A1(g8110A));
AND2_X1 U_g7930A (.ZN(g7930A),.A2(FE_OFN343_I5565A),.A1(g7621A));
AND3_X1 U_g8962A (.ZN(g8962A),.A3(g8828A),.A2(FE_OFN95_g2216A),.A1(g8089A));
AND2_X1 U_g10715A (.ZN(g10715A),.A2(g10584A),.A1(g2272A));
AND2_X1 U_g8659A (.ZN(g8659A),.A2(FE_OFN298_g3015A),.A1(g8269A));
AND2_X4 U_g3015A (.ZN(g3015A),.A2(I6260A),.A1(g2028A));
AND2_X1 U_g9643A (.ZN(g9643A),.A2(FE_OFN39_g9223A),.A1(g950A));
AND2_X4 U_g9205A (.ZN(g9205A),.A2(g8957A),.A1(FE_OFN276_g48A));
AND2_X1 U_g5538A (.ZN(g5538A),.A2(FE_OFN288_g4263A),.A1(g1669A));
AND2_X1 U_g4000A (.ZN(g4000A),.A2(g2774A),.A1(g1744A));
AND2_X1 U_g4126A (.ZN(g4126A),.A2(g3060A),.A1(FE_OFN253_g1786A));
AND2_X1 U_g4400A (.ZN(g4400A),.A2(FE_OFN137_g3829A),.A1(g4088A));
AND2_X1 U_g2794A (.ZN(g2794A),.A2(I5887A),.A1(I5886A));
AND2_X1 U_g4760A (.ZN(g4760A),.A2(FE_OFN307_g4010A),.A1(g486A));
AND2_X1 U_g6238A (.ZN(g6238A),.A2(FE_OFN289_g4679A),.A1(g572A));
AND2_X1 U_g10784A (.ZN(g10784A),.A2(g4467A),.A1(g10727A));
AND2_X1 U_g8174A (.ZN(g8174A),.A2(FE_OFN89_I11360A),.A1(g38A));
AND2_X1 U_g6332A (.ZN(g6332A),.A2(FE_OFN180_g5354A),.A1(g1374A));
AND2_X1 U_g5067A (.ZN(g5067A),.A2(g4811A),.A1(g305A));
AND2_X1 U_g5418A (.ZN(g5418A),.A2(FE_OFN357_g3521A),.A1(g1512A));
AND2_X1 U_g10297A (.ZN(g10297A),.A2(g10001A),.A1(FE_OFN79_g8700A));
AND2_X1 U_g6353A (.ZN(g6353A),.A2(FE_OFN320_g5361A),.A1(g299A));
AND2_X1 U_g11026A (.ZN(g11026A),.A2(FE_OFN14_g10702A),.A1(g386A));
AND2_X1 U_g11212A (.ZN(g11212A),.A2(FE_OFN279_g11157A),.A1(g944A));
AND2_X1 U_g6744A (.ZN(g6744A),.A2(FE_OFN218_g5557A),.A1(g4828A));
AND2_X1 U_g5493A (.ZN(g5493A),.A2(FE_OFN333_g4294A),.A1(g1923A));
AND2_X1 U_g10671A (.ZN(g10671A),.A2(g9473A),.A1(g10411A));
AND2_X1 U_g4383A (.ZN(g4383A),.A2(FE_OFN141_g3829A),.A1(g2517A));
AND2_X1 U_g5256A (.ZN(g5256A),.A2(g627A),.A1(g4297A));
AND2_X1 U_g4220A (.ZN(g4220A),.A2(g3539A),.A1(g105A));
AND2_X1 U_g8380A (.ZN(g8380A),.A2(FE_OFN333_g4294A),.A1(g8252A));
AND2_X1 U_g7071A (.ZN(g7071A),.A2(g6586A),.A1(g5030A));
AND2_X1 U_g4779A (.ZN(g4779A),.A2(FE_OFN307_g4010A),.A1(g501A));
AND2_X1 U_g9613A (.ZN(g9613A),.A2(FE_OFN46_g9125A),.A1(g1176A));
AND2_X1 U_g7705A (.ZN(g7705A),.A2(g4336A),.A1(g5935A));
AND2_X1 U_g9269A (.ZN(g9269A),.A2(FE_OFN266_g18A),.A1(g8933A));
AND2_X1 U_g5181A (.ZN(g5181A),.A2(g802A),.A1(g806A));
AND2_X1 U_g4977A (.ZN(g4977A),.A2(g4807A),.A1(g4567A));
AND2_X1 U_g7948A (.ZN(g7948A),.A2(g7497A),.A1(g70A));
AND2_X1 U_g11149A (.ZN(g11149A),.A2(FE_OFN278_g10927A),.A1(g324A));
AND2_X1 U_g9862A (.ZN(g9862A),.A2(g9778A),.A1(g1601A));
AND2_X1 U_g11387A (.ZN(g11387A),.A2(g3629A),.A1(g11077A));
AND2_X1 U_g7955A (.ZN(g7955A),.A2(g7516A),.A1(g76A));
AND2_X1 U_g4161A (.ZN(g4161A),.A2(g3060A),.A1(FE_OFN251_g1801A));
AND2_X1 U_g11148A (.ZN(g11148A),.A2(g10788A),.A1(g2321A));
AND2_X1 U_g9712A (.ZN(g9712A),.A2(FE_OFN70_g9490A),.A1(g1528A));
AND2_X1 U_g8931A (.ZN(g8931A),.A2(g8164A),.A1(g8642A));
AND2_X1 U_g11097A (.ZN(g11097A),.A2(g10883A),.A1(g378A));
AND3_X1 U_g5421A (.ZN(g5421A),.A3(g3819A),.A2(g109A),.A1(FE_OFN184_I7048A));
AND2_X1 U_g11104A (.ZN(g11104A),.A2(g10937A),.A1(g2963A));
AND2_X1 U_g5263A (.ZN(g5263A),.A2(FE_OFN335_g4737A),.A1(g709A));
AND2_X1 U_g6092A (.ZN(g6092A),.A2(FE_OFN273_g85A),.A1(g1059A));
AND2_X1 U_g4999A (.ZN(g4999A),.A2(FE_OFN154_g4640A),.A1(g1499A));
AND4_X1 U_I6338A (.ZN(I6338A),.A4(g2446A),.A3(g2451A),.A2(g2456A),.A1(g2475A));
AND3_X1 U_g7409A (.ZN(g7409A),.A3(g6858A),.A2(g632A),.A1(g4976A));
AND2_X1 U_g4103A (.ZN(g4103A),.A2(g3060A),.A1(FE_OFN247_g1771A));
AND4_X1 U_I6309A (.ZN(I6309A),.A4(g2475A),.A3(g2456A),.A2(g2451A),.A1(g2446A));
AND2_X1 U_g6580A (.ZN(g6580A),.A2(g5944A),.A1(FE_OFN251_g1801A));
AND2_X1 U_g5631A (.ZN(g5631A),.A2(FE_OFN291_g4880A),.A1(g1056A));
AND2_X1 U_g9414A (.ZN(g9414A),.A2(g9052A),.A1(g1730A));
AND2_X1 U_g9660A (.ZN(g9660A),.A2(FE_OFN45_g9125A),.A1(g1188A));
AND2_X1 U_g9946A (.ZN(g9946A),.A2(FE_OFN68_g9392A),.A1(g9926A));
AND2_X1 U_g5257A (.ZN(g5257A),.A2(FE_OFN335_g4737A),.A1(g691A));
AND2_X1 U_g4732A (.ZN(g4732A),.A2(FE_OFN300_g4002A),.A1(g391A));
AND2_X1 U_g3108A (.ZN(g3108A),.A2(I6331A),.A1(I6330A));
AND2_X1 U_g4753A (.ZN(g4753A),.A2(FE_OFN307_g4010A),.A1(g481A));
AND2_X1 U_g9903A (.ZN(g9903A),.A2(g9673A),.A1(g9885A));
AND2_X1 U_g10625A (.ZN(g10625A),.A2(FE_OFN369_g4525A),.A1(g10454A));
AND2_X1 U_g5605A (.ZN(g5605A),.A2(g704A),.A1(g4828A));
AND2_X1 U_g6623A (.ZN(g6623A),.A2(FE_OFN97_I8869A),.A1(g55A));
AND2_X1 U_g11228A (.ZN(g11228A),.A2(g11060A),.A1(g466A));
AND2_X1 U_g11011A (.ZN(g11011A),.A2(g10809A),.A1(g1968A));
AND2_X1 U_g6889A (.ZN(g6889A),.A2(FE_OFN213_g6003A),.A1(g1941A));
AND2_X1 U_g8040A (.ZN(g8040A),.A2(FE_OFN305_g5151A),.A1(g7523A));
AND2_X1 U_g7822A (.ZN(g7822A),.A2(FE_OFN209_g6863A),.A1(g1914A));
AND2_X1 U_g8123A (.ZN(g8123A),.A2(g7952A),.A1(g1918A));
AND2_X1 U_g11582A (.ZN(g11582A),.A2(g11539A),.A1(g1311A));
AND2_X1 U_g4316A (.ZN(g4316A),.A2(g3275A),.A1(g1965A));
AND2_X1 U_g10969A (.ZN(g10969A),.A2(g10809A),.A1(g3625A));
AND2_X1 U_g5041A (.ZN(g5041A),.A2(FE_OFN223_g4401A),.A1(g3983A));
AND2_X1 U_g9335A (.ZN(g9335A),.A2(FE_OFN275_g48A),.A1(g8975A));
AND2_X1 U_g9831A (.ZN(g9831A),.A2(FE_OFN34_g9785A),.A1(g9727A));
AND2_X1 U_g4565A (.ZN(g4565A),.A2(g4010A),.A1(g534A));
AND2_X1 U_g9422A (.ZN(g9422A),.A2(FE_OFN50_g9030A),.A1(g1750A));
AND2_X1 U_g8648A (.ZN(g8648A),.A2(g8511A),.A1(g4588A));
AND3_X1 U_g8875A (.ZN(g8875A),.A3(g8858A),.A2(FE_OFN92_g2216A),.A1(g8255A));
AND2_X1 U_g5168A (.ZN(g5168A),.A2(g4679A),.A1(g1512A));
AND2_X1 U_g7895A (.ZN(g7895A),.A2(FE_OFN334_g7045A),.A1(g7503A));
AND2_X1 U_g8655A (.ZN(g8655A),.A2(FE_OFN298_g3015A),.A1(g8267A));
AND2_X1 U_g4914A (.ZN(g4914A),.A2(FE_OFN290_g4880A),.A1(g1062A));
AND2_X1 U_g9947A (.ZN(g9947A),.A2(g9392A),.A1(g9927A));
AND2_X1 U_g5772A (.ZN(g5772A),.A2(FE_OFN321_g5261A),.A1(g1555A));
AND2_X1 U_g6838A (.ZN(g6838A),.A2(FE_OFN180_g5354A),.A1(g192A));
AND2_X1 U_g5531A (.ZN(g5531A),.A2(g4290A),.A1(g1666A));
AND2_X1 U_g6795A (.ZN(g6795A),.A2(g5878A),.A1(g5036A));
AND2_X1 U_g10503A (.ZN(g10503A),.A2(FE_OFN336_g1690A),.A1(g9995A));
AND2_X1 U_g8010A (.ZN(g8010A),.A2(g7438A),.A1(g7738A));
AND2_X1 U_g8410A (.ZN(g8410A),.A2(g8146A),.A1(g713A));
AND2_X1 U_g6231A (.ZN(g6231A),.A2(g5608A),.A1(g818A));
AND2_X1 U_g10581A (.ZN(g10581A),.A2(g9473A),.A1(g10336A));
AND2_X1 U_g10450A (.ZN(g10450A),.A2(FE_OFN235_g2024A),.A1(g10364A));
AND2_X1 U_g2804A (.ZN(g2804A),.A2(g1891A),.A1(g2132A));
AND2_X1 U_g3418A (.ZN(g3418A),.A2(FE_OFN352_g109A),.A1(g2379A));
AND2_X1 U_g9653A (.ZN(g9653A),.A2(FE_OFN45_g9125A),.A1(g1185A));
AND2_X1 U_g6205A (.ZN(g6205A),.A2(FE_OFN306_g5128A),.A1(g1515A));
AND2_X1 U_g10818A (.ZN(g10818A),.A2(FE_OFN204_g3664A),.A1(I16220A));
AND2_X1 U_g8172A (.ZN(g8172A),.A2(FE_OFN89_I11360A),.A1(g37A));
AND2_X1 U_g10496A (.ZN(g10496A),.A2(FE_OFN234_g2024A),.A1(g10429A));
AND2_X1 U_g5074A (.ZN(g5074A),.A2(g4608A),.A1(g1771A));
AND2_X1 U_g9869A (.ZN(g9869A),.A2(g9814A),.A1(g1558A));
AND2_X1 U_g9719A (.ZN(g9719A),.A2(g9490A),.A1(g1543A));
AND2_X1 U_g10741A (.ZN(g10741A),.A2(FE_OFN133_g3015A),.A1(g10635A));
AND2_X1 U_g3381A (.ZN(g3381A),.A2(g2756A),.A1(g940A));
AND2_X1 U_g5863A (.ZN(g5863A),.A2(g622A),.A1(g255A));
AND2_X1 U_g8693A (.ZN(g8693A),.A2(g8509A),.A1(g3738A));
AND2_X1 U_g5480A (.ZN(g5480A),.A2(FE_OFN366_g3521A),.A1(g554A));
AND2_X1 U_g4581A (.ZN(g4581A),.A2(g2047A),.A1(g3766A));
AND2_X1 U_g3685A (.ZN(g3685A),.A2(g2981A),.A1(FE_OFN238_g1781A));
AND2_X1 U_g5569A (.ZN(g5569A),.A2(g2338A),.A1(g4816A));
AND2_X1 U_g8555A (.ZN(g8555A),.A2(FE_OFN189_g7638A),.A1(g8409A));
AND2_X1 U_g3263A (.ZN(g3263A),.A2(g2328A),.A1(g2503A));
AND2_X1 U_g9364A (.ZN(g9364A),.A2(g9223A),.A1(g965A));
AND2_X1 U_g4784A (.ZN(g4784A),.A2(FE_OFN307_g4010A),.A1(g506A));
AND2_X4 U_g9454A (.ZN(g9454A),.A2(FE_OFN275_g48A),.A1(g8994A));
AND4_X1 U_I6331A (.ZN(I6331A),.A4(g2077A),.A3(g2074A),.A2(g2070A),.A1(g2060A));
AND2_X1 U_g11299A (.ZN(g11299A),.A2(g11243A),.A1(g4576A));
AND2_X1 U_g6983A (.ZN(g6983A),.A2(FE_OFN343_I5565A),.A1(g6592A));
AND2_X1 U_g7958A (.ZN(g7958A),.A2(FE_OFN198_g7697A),.A1(g736A));
AND2_X1 U_g4995A (.ZN(g4995A),.A2(FE_OFN153_g4640A),.A1(g1474A));
AND2_X1 U_g4079A (.ZN(g4079A),.A2(g2276A),.A1(FE_OFN237_g1806A));
AND2_X1 U_g2264A (.ZN(g2264A),.A2(g1766A),.A1(FE_OFN247_g1771A));
AND2_X1 U_g2160A (.ZN(g2160A),.A2(g746A),.A1(g745A));
AND2_X1 U_g3257A (.ZN(g3257A),.A2(g2496A),.A1(g378A));
AND2_X1 U_g3101A (.ZN(g3101A),.A2(I6310A),.A1(I6309A));
AND2_X1 U_g5000A (.ZN(g5000A),.A2(FE_OFN153_g4640A),.A1(g1470A));
AND2_X1 U_g3301A (.ZN(g3301A),.A2(g2544A),.A1(g1346A));
AND2_X1 U_g5126A (.ZN(g5126A),.A2(g4671A),.A1(g1104A));
AND4_X1 U_I5084A (.ZN(I5084A),.A4(g1478A),.A3(g1474A),.A2(g1470A),.A1(g1462A));
AND2_X1 U_g9412A (.ZN(g9412A),.A2(g9052A),.A1(g1727A));
AND2_X1 U_g9389A (.ZN(g9389A),.A2(FE_OFN47_g9151A),.A1(g1330A));
AND2_X1 U_g2379A (.ZN(g2379A),.A2(g743A),.A1(g744A));
AND2_X1 U_g10706A (.ZN(g10706A),.A2(FE_OFN345_g3015A),.A1(g10567A));
AND3_X1 U_I16145A (.ZN(I16145A),.A3(g10446A),.A2(g10447A),.A1(g10366A));
AND2_X1 U_g10597A (.ZN(g10597A),.A2(FE_OFN369_g4525A),.A1(g10533A));
AND3_X1 U_g8965A (.ZN(g8965A),.A3(g8849A),.A2(FE_OFN281_g2216A),.A1(g8110A));
AND2_X1 U_g5608A (.ZN(g5608A),.A2(g4831A),.A1(g814A));
AND2_X1 U_g5220A (.ZN(g5220A),.A2(g4776A),.A1(g1083A));
AND2_X1 U_g10624A (.ZN(g10624A),.A2(FE_OFN370_g4525A),.A1(g10494A));
AND2_X1 U_g10300A (.ZN(g10300A),.A2(g10019A),.A1(FE_OFN76_g8700A));
AND2_X1 U_g5023A (.ZN(g5023A),.A2(FE_OFN288_g4263A),.A1(g1071A));
AND2_X1 U_g4432A (.ZN(g4432A),.A2(g1975A),.A1(g3723A));
AND2_X1 U_g4053A (.ZN(g4053A),.A2(FE_OFN224_g2276A),.A1(FE_OFN253_g1786A));
AND2_X1 U_g8050A (.ZN(g8050A),.A2(FE_OFN177_g5919A),.A1(g7596A));
AND2_X1 U_g5588A (.ZN(g5588A),.A2(FE_OFN367_g3521A),.A1(g1639A));
AND3_X1 U_g6679A (.ZN(g6679A),.A3(g109A),.A2(g6074A),.A1(FE_OFN184_I7048A));
AND2_X1 U_g9963A (.ZN(g9963A),.A2(FE_OFN280_g9536A),.A1(g9953A));
AND2_X1 U_g3772A (.ZN(g3772A),.A2(g3089A),.A1(g2542A));
AND2_X1 U_g5051A (.ZN(g5051A),.A2(g2506A),.A1(g4432A));
AND2_X1 U_g6831A (.ZN(g6831A),.A2(FE_OFN179_g5354A),.A1(g207A));
AND2_X1 U_g2981A (.ZN(g2981A),.A2(g2264A),.A1(FE_OFN236_g1776A));
AND2_X1 U_g8724A (.ZN(g8724A),.A2(g7910A),.A1(g8214A));
AND2_X1 U_g4157A (.ZN(g4157A),.A2(g3060A),.A1(FE_OFN239_g1796A));
AND2_X1 U_g9707A (.ZN(g9707A),.A2(g9474A),.A1(g1583A));
AND3_X1 U_g8878A (.ZN(g8878A),.A3(FE_OFN73_g8858A),.A2(FE_OFN93_g2216A),.A1(g8099A));
AND2_X1 U_g2132A (.ZN(g2132A),.A2(g1882A),.A1(g1872A));
AND2_X1 U_g10763A (.ZN(g10763A),.A2(FE_OFN345_g3015A),.A1(g10639A));
AND3_X1 U_g8289A (.ZN(g8289A),.A3(g2216A),.A2(g8109A),.A1(g6777A));
AND2_X1 U_g7898A (.ZN(g7898A),.A2(g7045A),.A1(g7511A));
AND2_X1 U_g11271A (.ZN(g11271A),.A2(g11203A),.A1(g4753A));
AND2_X1 U_g11461A (.ZN(g11461A),.A2(FE_OFN100_g4421A),.A1(g11225A));
AND2_X1 U_g5732A (.ZN(g5732A),.A2(FE_OFN353_g5117A),.A1(g1604A));
AND2_X1 U_g11145A (.ZN(g11145A),.A2(FE_OFN278_g10927A),.A1(g315A));
AND2_X1 U_g11031A (.ZN(g11031A),.A2(FE_OFN14_g10702A),.A1(g411A));
AND2_X1 U_g9865A (.ZN(g9865A),.A2(g9773A),.A1(g1607A));
AND2_X1 U_g5944A (.ZN(g5944A),.A2(g5233A),.A1(g1796A));
AND2_X1 U_g9715A (.ZN(g9715A),.A2(FE_OFN70_g9490A),.A1(g1531A));
AND2_X1 U_g9604A (.ZN(g9604A),.A2(FE_OFN51_g9111A),.A1(g1194A));
AND2_X1 U_g8799A (.ZN(g8799A),.A2(FE_OFN331_g8696A),.A1(g8647A));
AND2_X1 U_g11198A (.ZN(g11198A),.A2(FE_OFN15_g10702A),.A1(g4778A));
AND2_X1 U_g6873A (.ZN(g6873A),.A2(g6557A),.A1(g3263A));
AND2_X1 U_g6632A (.ZN(g6632A),.A2(FE_OFN283_I8869A),.A1(g61A));
AND2_X1 U_g6095A (.ZN(g6095A),.A2(FE_OFN273_g85A),.A1(g1062A));
AND2_X1 U_g3863A (.ZN(g3863A),.A2(g1696A),.A1(g1703A));
AND2_X1 U_g9833A (.ZN(g9833A),.A2(FE_OFN34_g9785A),.A1(g9729A));
AND2_X1 U_g6653A (.ZN(g6653A),.A2(I8869A),.A1(g70A));
AND2_X1 U_g6102A (.ZN(g6102A),.A2(FE_OFN273_g85A),.A1(g1038A));
AND2_X1 U_g7819A (.ZN(g7819A),.A2(FE_OFN206_g6863A),.A1(g1887A));
AND2_X1 U_g11393A (.ZN(g11393A),.A2(g7914A),.A1(g11280A));
AND2_X1 U_g2511A (.ZN(g2511A),.A2(g456A),.A1(FE_OFN254_g461A));
AND2_X1 U_g7088A (.ZN(g7088A),.A2(g6432A),.A1(g2331A));
AND2_X1 U_g9584A (.ZN(g9584A),.A2(FE_OFN53_g9173A),.A1(g1341A));
AND2_X1 U_g9896A (.ZN(g9896A),.A2(FE_OFN60_g9624A),.A1(g9696A));
AND3_X1 U_g8209A (.ZN(g8209A),.A3(g7622A),.A2(g3068A),.A1(g4094A));
AND2_X1 U_g6752A (.ZN(g6752A),.A2(g2343A),.A1(g6187A));
AND2_X1 U_g4778A (.ZN(g4778A),.A2(g4002A),.A1(g421A));
AND2_X1 U_g11161A (.ZN(g11161A),.A2(g10937A),.A1(g1969A));
AND2_X1 U_g9268A (.ZN(g9268A),.A2(g8947A),.A1(g6109A));
AND2_X1 U_g5681A (.ZN(g5681A),.A2(FE_OFN365_g5361A),.A1(g135A));
AND2_X1 U_g7951A (.ZN(g7951A),.A2(g7505A),.A1(g73A));
AND2_X1 U_g9419A (.ZN(g9419A),.A2(FE_OFN50_g9030A),.A1(g1744A));
AND2_X1 U_g10268A (.ZN(g10268A),.A2(FE_OFN267_g109A),.A1(I15287A));
AND2_X1 U_g5533A (.ZN(g5533A),.A2(g4292A),.A1(g1724A));
AND2_X4 U_g9052A (.ZN(g9052A),.A2(FE_OFN276_g48A),.A1(g8936A));
AND2_X1 U_g6786A (.ZN(g6786A),.A2(g5919A),.A1(g178A));
AND2_X1 U_g10670A (.ZN(g10670A),.A2(g9097A),.A1(g10396A));
AND2_X1 U_g11087A (.ZN(g11087A),.A2(FE_OFN4_g10950A),.A1(g829A));
AND2_X1 U_g4949A (.ZN(g4949A),.A2(g4449A),.A1(I5815A));
AND2_X1 U_g6364A (.ZN(g6364A),.A2(FE_OFN346_g4381A),.A1(g5851A));
AND2_X1 U_g7825A (.ZN(g7825A),.A2(FE_OFN206_g6863A),.A1(g1941A));
AND2_X1 U_g4998A (.ZN(g4998A),.A2(FE_OFN303_g4678A),.A1(g1304A));
AND2_X1 U_g10667A (.ZN(g10667A),.A2(g9424A),.A1(g10405A));
AND2_X1 U_g7136A (.ZN(g7136A),.A2(g6718A),.A1(g5190A));
AND2_X1 U_g6532A (.ZN(g6532A),.A2(FE_OFN282_g6165A),.A1(g339A));
AND2_X1 U_g9385A (.ZN(g9385A),.A2(FE_OFN48_g9151A),.A1(g1324A));
AND4_X1 U_I5690A (.ZN(I5690A),.A4(g1448A),.A3(g1444A),.A2(g1440A),.A1(g1436A));
AND2_X1 U_g4484A (.ZN(g4484A),.A2(FE_OFN302_g3913A),.A1(g1137A));
AND2_X1 U_g9897A (.ZN(g9897A),.A2(FE_OFN60_g9624A),.A1(g9699A));
AND2_X1 U_g9425A (.ZN(g9425A),.A2(FE_OFN49_g9030A),.A1(g1753A));
AND2_X1 U_g3383A (.ZN(g3383A),.A2(FE_OFN324_g18A),.A1(g186A));
AND2_X1 U_g5601A (.ZN(g5601A),.A2(g4880A),.A1(g1035A));
AND2_X1 U_g7943A (.ZN(g7943A),.A2(g7467A),.A1(g64A));
AND2_X1 U_g11171A (.ZN(g11171A),.A2(FE_OFN21_g10702A),.A1(g481A));
AND2_X1 U_g3423A (.ZN(g3423A),.A2(I6631A),.A1(I6630A));
AND2_X1 U_g7230A (.ZN(g7230A),.A2(g6447A),.A1(g6064A));
AND2_X1 U_g4952A (.ZN(g4952A),.A2(FE_OFN299_g4457A),.A1(g1648A));
AND2_X1 U_g6787A (.ZN(g6787A),.A2(FE_OFN319_g5361A),.A1(g266A));
AND3_X1 U_g8968A (.ZN(g8968A),.A3(g8849A),.A2(FE_OFN281_g2216A),.A1(g8089A));
AND2_X1 U_g10306A (.ZN(g10306A),.A2(g9082A),.A1(g10007A));
AND2_X1 U_g9331A (.ZN(g9331A),.A2(FE_OFN275_g48A),.A1(g8972A));
AND2_X1 U_g11459A (.ZN(g11459A),.A2(FE_OFN100_g4421A),.A1(g11221A));
AND2_X1 U_g4561A (.ZN(g4561A),.A2(g4010A),.A1(g538A));
AND2_X1 U_g11425A (.ZN(g11425A),.A2(g10629A),.A1(I16982A));
AND2_X1 U_g11458A (.ZN(g11458A),.A2(FE_OFN99_g4421A),.A1(g11219A));
AND2_X1 U_g5739A (.ZN(g5739A),.A2(FE_OFN315_g5117A),.A1(g1607A));
AND2_X1 U_g7496A (.ZN(g7496A),.A2(g64A),.A1(FE_OFN83_g2176A));
AND2_X1 U_g4986A (.ZN(g4986A),.A2(FE_OFN146_g4682A),.A1(g1411A));
AND2_X1 U_g11010A (.ZN(g11010A),.A2(FE_OFN18_g10702A),.A1(g5187A));
AND2_X1 U_g3999A (.ZN(g3999A),.A2(g2777A),.A1(g1741A));
AND2_X1 U_g8175A (.ZN(g8175A),.A2(FE_OFN89_I11360A),.A1(g39A));
AND2_X1 U_g8722A (.ZN(g8722A),.A2(g7908A),.A1(g8210A));
AND2_X1 U_g4764A (.ZN(g4764A),.A2(FE_OFN300_g4002A),.A1(g411A));
AND2_X1 U_g7137A (.ZN(g7137A),.A2(g6354A),.A1(g5590A));
AND2_X1 U_g7891A (.ZN(g7891A),.A2(FE_OFN334_g7045A),.A1(g7471A));
AND2_X1 U_g8651A (.ZN(g8651A),.A2(FE_OFN348_g3015A),.A1(g8261A));
AND2_X1 U_g5479A (.ZN(g5479A),.A2(g4243A),.A1(g1845A));
AND2_X1 U_g11599A (.ZN(g11599A),.A2(g11575A),.A1(g1341A));
AND2_X1 U_g6684A (.ZN(g6684A),.A2(g5836A),.A1(g91A));
AND2_X1 U_g6745A (.ZN(g6745A),.A2(FE_OFN218_g5557A),.A1(g5605A));
AND2_X1 U_g6639A (.ZN(g6639A),.A2(FE_OFN282_g6165A),.A1(g357A));
AND2_X1 U_g10937A (.ZN(g10937A),.A2(FE_OFN13_g10702A),.A1(g4822A));
AND2_X1 U_g3696A (.ZN(g3696A),.A2(FE_OFN364_g3015A),.A1(g1713A));
AND2_X1 U_g4503A (.ZN(g4503A),.A2(g3943A),.A1(g654A));
AND2_X1 U_g6791A (.ZN(g6791A),.A2(FE_OFN319_g5361A),.A1(g269A));
AND2_X1 U_g5190A (.ZN(g5190A),.A2(g4678A),.A1(g1245A));
AND2_X1 U_g5390A (.ZN(g5390A),.A2(g4671A),.A1(g1101A));
AND2_X1 U_g8384A (.ZN(g8384A),.A2(FE_OFN325_g18A),.A1(g8180A));
AND2_X1 U_g4224A (.ZN(g4224A),.A2(FE_OFN132_g3015A),.A1(g1092A));
AND2_X1 U_g5501A (.ZN(g5501A),.A2(g4273A),.A1(g1672A));
AND2_X4 U_g9173A (.ZN(g9173A),.A2(FE_OFN276_g48A),.A1(g8968A));
AND2_X1 U_g6759A (.ZN(g6759A),.A2(g5919A),.A1(g148A));
AND2_X1 U_g8838A (.ZN(g8838A),.A2(FE_OFN328_g8709A),.A1(g8602A));
AND2_X1 U_g8024A (.ZN(g8024A),.A2(FE_OFN322_g4449A),.A1(g6577A));
AND2_X1 U_g10666A (.ZN(g10666A),.A2(g9424A),.A1(g10402A));
AND2_X1 U_g11158A (.ZN(g11158A),.A2(FE_OFN278_g10927A),.A1(g309A));
AND2_X1 U_g9602A (.ZN(g9602A),.A2(g9010A),.A1(g932A));
AND2_X1 U_g5704A (.ZN(g5704A),.A2(FE_OFN164_g5361A),.A1(g143A));
AND2_X1 U_g4617A (.ZN(g4617A),.A2(g3879A),.A1(g3275A));
AND2_X2 U_g11561A (.ZN(g11561A),.A2(FE_OFN364_g3015A),.A1(g11492A));
AND2_X1 U_g9868A (.ZN(g9868A),.A2(g9814A),.A1(g1555A));
AND2_X1 U_g11295A (.ZN(g11295A),.A2(g11239A),.A1(g4554A));
AND2_X1 U_g11144A (.ZN(g11144A),.A2(FE_OFN10_g10702A),.A1(g305A));
AND2_X1 U_g9718A (.ZN(g9718A),.A2(FE_OFN70_g9490A),.A1(g1540A));
AND2_X1 U_g3434A (.ZN(g3434A),.A2(g2355A),.A1(g237A));
AND2_X1 U_g4987A (.ZN(g4987A),.A2(FE_OFN147_g4682A),.A1(g1440A));
AND2_X1 U_g4771A (.ZN(g4771A),.A2(FE_OFN307_g4010A),.A1(g496A));
AND2_X1 U_g5250A (.ZN(g5250A),.A2(g4678A),.A1(g1270A));
AND2_X1 U_g6098A (.ZN(g6098A),.A2(FE_OFN273_g85A),.A1(g1065A));
AND2_X1 U_g9582A (.ZN(g9582A),.A2(FE_OFN53_g9173A),.A1(g2725A));
AND2_X1 U_g6833A (.ZN(g6833A),.A2(FE_OFN178_g5354A),.A1(g186A));
AND2_X1 U_g3533A (.ZN(g3533A),.A2(g2892A),.A1(g1981A));
AND2_X1 U_g4892A (.ZN(g4892A),.A2(g4739A),.A1(g632A));
AND2_X1 U_g8104A (.ZN(g8104A),.A2(g7852A),.A1(g5493A));
AND2_X1 U_g9415A (.ZN(g9415A),.A2(FE_OFN54_g9052A),.A1(g1733A));
AND2_X1 U_g8499A (.ZN(g8499A),.A2(g4737A),.A1(g8377A));
AND2_X1 U_g9664A (.ZN(g9664A),.A2(FE_OFN46_g9125A),.A1(g1191A));
AND2_X1 U_g9721A (.ZN(g9721A),.A2(FE_OFN359_g18A),.A1(g9413A));
AND2_X1 U_g6162A (.ZN(g6162A),.A2(g5200A),.A1(g3584A));
AND2_X1 U_g4991A (.ZN(g4991A),.A2(FE_OFN154_g4640A),.A1(g1508A));
AND2_X1 U_g6362A (.ZN(g6362A),.A2(FE_OFN346_g4381A),.A1(g5846A));
AND4_X1 U_I6631A (.ZN(I6631A),.A4(FE_OFN237_g1806A),.A3(FE_OFN251_g1801A),.A2(FE_OFN239_g1796A),.A1(FE_OFN252_g1791A));
AND2_X1 U_g10685A (.ZN(g10685A),.A2(FE_OFN136_g3863A),.A1(g10383A));
AND2_X1 U_g4340A (.ZN(g4340A),.A2(FE_OFN351_g3913A),.A1(g1153A));
AND2_X1 U_g11023A (.ZN(g11023A),.A2(g10702A),.A1(g440A));
AND2_X1 U_g8044A (.ZN(g8044A),.A2(FE_OFN177_g5919A),.A1(g7598A));
AND2_X1 U_g11224A (.ZN(g11224A),.A2(g11157A),.A1(g968A));
AND2_X1 U_g11571A (.ZN(g11571A),.A2(g11561A),.A1(g2018A));
AND2_X1 U_g4959A (.ZN(g4959A),.A2(FE_OFN147_g4682A),.A1(g1520A));
AND2_X1 U_g10334A (.ZN(g10334A),.A2(FE_OFN267_g109A),.A1(I15365A));
AND2_X1 U_g5626A (.ZN(g5626A),.A2(FE_OFN367_g3521A),.A1(g1633A));
AND2_X1 U_g9940A (.ZN(g9940A),.A2(FE_OFN67_g9367A),.A1(g9920A));
AND2_X1 U_g4876A (.ZN(g4876A),.A2(FE_OFN132_g3015A),.A1(g1086A));
AND2_X1 U_g6728A (.ZN(g6728A),.A2(FE_OFN310_g4336A),.A1(g4482A));
AND2_X1 U_g6730A (.ZN(g6730A),.A2(g5013A),.A1(g1872A));
AND2_X1 U_g9689A (.ZN(g9689A),.A2(FE_OFN59_g9432A),.A1(g263A));
AND2_X1 U_g10762A (.ZN(g10762A),.A2(FE_OFN131_g3015A),.A1(g10635A));
AND2_X1 U_g6070A (.ZN(g6070A),.A2(FE_OFN273_g85A),.A1(g1050A));
AND2_X1 U_g9428A (.ZN(g9428A),.A2(FE_OFN50_g9030A),.A1(g1756A));
AND2_X4 U_g9030A (.ZN(g9030A),.A2(FE_OFN276_g48A),.A1(g8935A));
AND2_X1 U_g9430A (.ZN(g9430A),.A2(FE_OFN49_g9030A),.A1(g1759A));
AND2_X1 U_g8927A (.ZN(g8927A),.A2(g8642A),.A1(g2216A));
AND2_X1 U_g7068A (.ZN(g7068A),.A2(g6586A),.A1(g5024A));
AND2_X1 U_g8014A (.ZN(g8014A),.A2(g7438A),.A1(g7740A));
AND2_X1 U_g11392A (.ZN(g11392A),.A2(g7914A),.A1(g11278A));
AND2_X1 U_g5782A (.ZN(g5782A),.A2(g5222A),.A1(g1558A));
AND2_X1 U_g4824A (.ZN(g4824A),.A2(g4099A),.A1(g774A));
AND2_X1 U_g6331A (.ZN(g6331A),.A2(FE_OFN180_g5354A),.A1(g201A));
AND2_X1 U_g4236A (.ZN(g4236A),.A2(FE_OFN132_g3015A),.A1(g1098A));
AND2_X1 U_g11559A (.ZN(g11559A),.A2(FE_OFN27_g11519A),.A1(FE_OFN251_g1801A));
AND2_X1 U_g9609A (.ZN(g9609A),.A2(FE_OFN42_g9205A),.A1(g907A));
AND2_X1 U_g11558A (.ZN(g11558A),.A2(FE_OFN27_g11519A),.A1(FE_OFN239_g1796A));
AND2_X1 U_g6087A (.ZN(g6087A),.A2(FE_OFN271_g85A),.A1(g1056A));
AND2_X1 U_g5526A (.ZN(g5526A),.A2(g4294A),.A1(g1950A));
AND2_X1 U_g10751A (.ZN(g10751A),.A2(FE_OFN133_g3015A),.A1(g10646A));
AND2_X1 U_g10772A (.ZN(g10772A),.A2(FE_OFN345_g3015A),.A1(g10655A));
AND2_X1 U_g8135A (.ZN(g8135A),.A2(g7883A),.A1(g1945A));
AND2_X1 U_g11544A (.ZN(g11544A),.A2(g10584A),.A1(g11515A));
AND2_X1 U_g5084A (.ZN(g5084A),.A2(FE_OFN299_g4457A),.A1(g1776A));
AND2_X1 U_g8382A (.ZN(g8382A),.A2(FE_OFN196_g7697A),.A1(g5248A));
AND2_X1 U_g10230A (.ZN(g10230A),.A2(g9968A),.A1(g8700A));
AND2_X1 U_g5484A (.ZN(g5484A),.A2(FE_OFN333_g4294A),.A1(g1896A));
AND2_X1 U_g7241A (.ZN(g7241A),.A2(g5557A),.A1(g6772A));
AND2_X1 U_g3942A (.ZN(g3942A),.A2(FE_OFN260_g18A),.A1(g219A));
AND2_X1 U_g10638A (.ZN(g10638A),.A2(g3829A),.A1(g10383A));
AND2_X1 U_g4064A (.ZN(g4064A),.A2(g2774A),.A1(g1759A));
AND2_X1 U_g9365A (.ZN(g9365A),.A2(FE_OFN48_g9151A),.A1(g1321A));
AND2_X1 U_g9861A (.ZN(g9861A),.A2(g9579A),.A1(g9738A));
AND2_X1 U_g11255A (.ZN(g11255A),.A2(g11060A),.A1(g456A));
AND2_X1 U_g11189A (.ZN(g11189A),.A2(FE_OFN15_g10702A),.A1(g4736A));
AND2_X1 U_g10510A (.ZN(g10510A),.A2(FE_OFN336_g1690A),.A1(g10019A));
AND3_X1 U_g8947A (.ZN(g8947A),.A3(g8828A),.A2(FE_OFN92_g2216A),.A1(g8056A));
AND2_X1 U_g2917A (.ZN(g2917A),.A2(g1657A),.A1(g2424A));
AND2_X2 U_g5919A (.ZN(g5919A),.A2(FE_OFN269_g109A),.A1(I7048A));
AND2_X1 U_g11188A (.ZN(g11188A),.A2(FE_OFN15_g10702A),.A1(g4732A));
AND2_X1 U_g9846A (.ZN(g9846A),.A2(g9764A),.A1(g287A));
AND2_X1 U_g7818A (.ZN(g7818A),.A2(FE_OFN206_g6863A),.A1(g1878A));
AND2_X1 U_g11460A (.ZN(g11460A),.A2(FE_OFN99_g4421A),.A1(g11223A));
AND2_X1 U_g5276A (.ZN(g5276A),.A2(FE_OFN335_g4737A),.A1(g736A));
AND2_X1 U_g11030A (.ZN(g11030A),.A2(FE_OFN17_g10702A),.A1(g406A));
AND2_X1 U_g11093A (.ZN(g11093A),.A2(FE_OFN4_g10950A),.A1(g841A));
AND2_X1 U_g7893A (.ZN(g7893A),.A2(FE_OFN334_g7045A),.A1(g7478A));
AND2_X1 U_g8653A (.ZN(g8653A),.A2(FE_OFN348_g3015A),.A1(g8265A));
AND2_X1 U_g10442A (.ZN(g10442A),.A2(FE_OFN245_g1690A),.A1(g9968A));
AND2_X1 U_g6535A (.ZN(g6535A),.A2(g6165A),.A1(g345A));
AND2_X1 U_g8102A (.ZN(g8102A),.A2(g7852A),.A1(g5485A));
AND4_X1 U_I5085A (.ZN(I5085A),.A4(g1508A),.A3(g1504A),.A2(g1494A),.A1(g1490A));
AND2_X1 U_g5004A (.ZN(g5004A),.A2(FE_OFN303_g4678A),.A1(g1296A));
AND2_X1 U_g3912A (.ZN(g3912A),.A2(FE_OFN359_g18A),.A1(g207A));
AND2_X1 U_g7186A (.ZN(g7186A),.A2(g6403A),.A1(g2503A));
AND2_X1 U_g4489A (.ZN(g4489A),.A2(FE_OFN103_g3586A),.A1(g348A));
AND2_X1 U_g9662A (.ZN(g9662A),.A2(g9292A),.A1(g123A));
AND2_X1 U_g9418A (.ZN(g9418A),.A2(FE_OFN56_g9052A),.A1(g1741A));
AND2_X1 U_g11218A (.ZN(g11218A),.A2(FE_OFN279_g11157A),.A1(g959A));
AND2_X1 U_g4471A (.ZN(g4471A),.A2(FE_OFN302_g3913A),.A1(g1121A));
AND2_X1 U_g10746A (.ZN(g10746A),.A2(FE_OFN364_g3015A),.A1(g10643A));
AND2_X1 U_g7125A (.ZN(g7125A),.A2(g5763A),.A1(g1212A));
AND2_X1 U_g7821A (.ZN(g7821A),.A2(FE_OFN209_g6863A),.A1(g1905A));
AND2_X1 U_g6246A (.ZN(g6246A),.A2(FE_OFN164_g5361A),.A1(g178A));
AND2_X1 U_g9256A (.ZN(g9256A),.A2(g8963A),.A1(g6109A));
AND2_X1 U_g8042A (.ZN(g8042A),.A2(FE_OFN305_g5151A),.A1(g7533A));
AND2_X1 U_g10237A (.ZN(g10237A),.A2(g9082A),.A1(g9968A));
AND2_X1 U_g7939A (.ZN(g7939A),.A2(g7460A),.A1(g61A));
AND2_X1 U_g8786A (.ZN(g8786A),.A2(FE_OFN331_g8696A),.A1(g8638A));
AND2_X1 U_g10684A (.ZN(g10684A),.A2(FE_OFN136_g3863A),.A1(g10382A));
AND2_X1 U_g11455A (.ZN(g11455A),.A2(FE_OFN99_g4421A),.A1(g11233A));
AND2_X1 U_g8364A (.ZN(g8364A),.A2(g8146A),.A1(g658A));
AND3_X1 U_g2990A (.ZN(g2990A),.A3(g1814A),.A2(g2557A),.A1(g2061A));
AND2_X1 U_g9847A (.ZN(g9847A),.A2(FE_OFN57_g9432A),.A1(g290A));
AND2_X1 U_g8054A (.ZN(g8054A),.A2(FE_OFN177_g5919A),.A1(g7584A));
AND2_X1 U_g5617A (.ZN(g5617A),.A2(FE_OFN290_g4880A),.A1(g1050A));
AND2_X1 U_g6502A (.ZN(g6502A),.A2(FE_OFN363_I5565A),.A1(g5981A));
AND2_X1 U_g5789A (.ZN(g5789A),.A2(FE_OFN321_g5261A),.A1(g1561A));
AND2_X1 U_g4009A (.ZN(g4009A),.A2(g2774A),.A1(g1747A));
AND2_X1 U_g11277A (.ZN(g11277A),.A2(g11199A),.A1(g4779A));
AND2_X1 U_g6940A (.ZN(g6940A),.A2(g1945A),.A1(g6472A));
AND2_X1 U_g7061A (.ZN(g7061A),.A2(g6760A),.A1(g790A));
AND2_X1 U_g11595A (.ZN(g11595A),.A2(g11575A),.A1(g1336A));
AND2_X1 U_g5771A (.ZN(g5771A),.A2(FE_OFN321_g5261A),.A1(g1534A));
AND2_X1 U_g8553A (.ZN(g8553A),.A2(FE_OFN330_g7638A),.A1(g8405A));
AND2_X1 U_g4836A (.ZN(g4836A),.A2(g3943A),.A1(g643A));
AND2_X1 U_g5547A (.ZN(g5547A),.A2(g4292A),.A1(g1733A));
AND2_X1 U_g6216A (.ZN(g6216A),.A2(FE_OFN306_g5128A),.A1(g1407A));
AND2_X1 U_g4967A (.ZN(g4967A),.A2(FE_OFN146_g4682A),.A1(g1515A));
AND2_X1 U_g6671A (.ZN(g6671A),.A2(FE_OFN282_g6165A),.A1(g342A));
AND2_X1 U_g7200A (.ZN(g7200A),.A2(g6447A),.A1(g3098A));
AND2_X1 U_g3661A (.ZN(g3661A),.A2(g3257A),.A1(g382A));
AND2_X1 U_g7046A (.ZN(g7046A),.A2(g6702A),.A1(g4998A));
AND2_X1 U_g4229A (.ZN(g4229A),.A2(g4673A),.A1(g999A));
AND2_X1 U_g8389A (.ZN(g8389A),.A2(g8220A),.A1(g5263A));
AND2_X1 U_g6430A (.ZN(g6430A),.A2(FE_OFN217_g5013A),.A1(g5044A));
AND2_X1 U_g4993A (.ZN(g4993A),.A2(FE_OFN147_g4682A),.A1(g1448A));
AND2_X1 U_g6247A (.ZN(g6247A),.A2(FE_OFN365_g5361A),.A1(g127A));
AND2_X1 U_g9257A (.ZN(g9257A),.A2(g8964A),.A1(g6109A));
AND2_X1 U_g11170A (.ZN(g11170A),.A2(FE_OFN8_g10702A),.A1(g525A));
AND2_X1 U_g7145A (.ZN(g7145A),.A2(g6718A),.A1(g5250A));
AND2_X1 U_g5738A (.ZN(g5738A),.A2(FE_OFN353_g5117A),.A1(g1586A));
AND2_X1 U_g6826A (.ZN(g6826A),.A2(g5354A),.A1(g225A));
AND2_X1 U_g7191A (.ZN(g7191A),.A2(FE_OFN310_g4336A),.A1(g5219A));
AND2_X1 U_g3998A (.ZN(g3998A),.A2(g2276A),.A1(g2677A));
AND2_X1 U_g6741A (.ZN(g6741A),.A2(FE_OFN219_g5557A),.A1(g3284A));
AND2_X1 U_g5478A (.ZN(g5478A),.A2(FE_OFN333_g4294A),.A1(g1905A));
AND2_X1 U_g11167A (.ZN(g11167A),.A2(FE_OFN8_g10702A),.A1(g538A));
AND2_X1 U_g11194A (.ZN(g11194A),.A2(g10927A),.A1(g4764A));
AND2_X1 U_g11589A (.ZN(g11589A),.A2(g11539A),.A1(g1333A));
AND2_X1 U_g6638A (.ZN(g6638A),.A2(FE_OFN283_I8869A),.A1(g64A));
AND2_X2 U_g4921A (.ZN(g4921A),.A2(g4431A),.A1(g627A));
AND2_X1 U_g7536A (.ZN(g7536A),.A2(g76A),.A1(FE_OFN83_g2176A));
AND2_X1 U_g9585A (.ZN(g9585A),.A2(g8995A),.A1(g889A));
AND2_X1 U_g2957A (.ZN(g2957A),.A2(g1663A),.A1(g2424A));
AND2_X1 U_g11588A (.ZN(g11588A),.A2(g11547A),.A1(g1330A));
AND2_X1 U_g5690A (.ZN(g5690A),.A2(FE_OFN353_g5117A),.A1(g1567A));
AND2_X1 U_g6883A (.ZN(g6883A),.A2(FE_OFN213_g6003A),.A1(g1923A));
AND2_X1 U_g4837A (.ZN(g4837A),.A2(FE_OFN297_g3015A),.A1(g1068A));
AND3_X1 U_g8963A (.ZN(g8963A),.A3(g8849A),.A2(FE_OFN92_g2216A),.A1(g8056A));
AND2_X1 U_g8791A (.ZN(g8791A),.A2(FE_OFN331_g8696A),.A1(g8641A));
AND2_X1 U_g6217A (.ZN(g6217A),.A2(FE_OFN291_g4880A),.A1(g563A));
AND4_X1 U_I6316A (.ZN(I6316A),.A4(g2395A),.A3(g2381A),.A2(g2087A),.A1(g2082A));
AND2_X1 U_g11022A (.ZN(g11022A),.A2(g10702A),.A1(g444A));
AND2_X1 U_g5915A (.ZN(g5915A),.A2(g4977A),.A1(g4168A));
AND2_X1 U_g4788A (.ZN(g4788A),.A2(FE_OFN307_g4010A),.A1(g511A));
AND2_X1 U_g5110A (.ZN(g5110A),.A2(FE_OFN299_g4457A),.A1(FE_OFN237_g1806A));
AND2_X1 U_g11254A (.ZN(g11254A),.A2(g11083A),.A1(g986A));
AND2_X1 U_g6827A (.ZN(g6827A),.A2(FE_OFN178_g5354A),.A1(g219A));
AND3_X1 U_g8957A (.ZN(g8957A),.A3(g8828A),.A2(FE_OFN281_g2216A),.A1(g8081A));
AND2_X1 U_g6333A (.ZN(g6333A),.A2(FE_OFN180_g5354A),.A1(g197A));
AND2_X1 U_g8049A (.ZN(g8049A),.A2(FE_OFN177_g5919A),.A1(g7567A));
AND2_X1 U_g4392A (.ZN(g4392A),.A2(FE_OFN137_g3829A),.A1(g3273A));
AND2_X1 U_g9856A (.ZN(g9856A),.A2(g9773A),.A1(g1592A));
AND2_X1 U_g9411A (.ZN(g9411A),.A2(g9052A),.A1(g1724A));
AND2_X1 U_g5002A (.ZN(g5002A),.A2(FE_OFN154_g4640A),.A1(g1494A));
AND2_X1 U_g11101A (.ZN(g11101A),.A2(FE_OFN4_g10950A),.A1(g857A));
AND2_X1 U_g11177A (.ZN(g11177A),.A2(FE_OFN20_g10702A),.A1(g511A));
AND2_X1 U_g11560A (.ZN(g11560A),.A2(FE_OFN27_g11519A),.A1(g1806A));
AND2_X1 U_g8098A (.ZN(g8098A),.A2(g7852A),.A1(g5478A));
AND2_X1 U_g3970A (.ZN(g3970A),.A2(FE_OFN260_g18A),.A1(g225A));
AND2_X1 U_g4941A (.ZN(g4941A),.A2(FE_OFN290_g4880A),.A1(g1038A));
AND2_X1 U_g10453A (.ZN(g10453A),.A2(FE_OFN234_g2024A),.A1(g10437A));
AND2_X1 U_g5877A (.ZN(g5877A),.A2(g639A),.A1(g4921A));
AND2_X1 U_g6662A (.ZN(g6662A),.A2(FE_OFN282_g6165A),.A1(g366A));
AND2_X1 U_g7935A (.ZN(g7935A),.A2(g7454A),.A1(g58A));
AND2_X1 U_g6067A (.ZN(g6067A),.A2(g85A),.A1(g1047A));
AND4_X1 U_I6317A (.ZN(I6317A),.A4(g2438A),.A3(g2434A),.A2(g2420A),.A1(g2406A));
AND2_X1 U_g9863A (.ZN(g9863A),.A2(FE_OFN56_g9052A),.A1(g9740A));
AND4_X1 U_I5886A (.ZN(I5886A),.A4(g2254A),.A3(g2249A),.A2(g170A),.A1(g174A));
AND2_X1 U_g6994A (.ZN(g6994A),.A2(FE_OFN141_g3829A),.A1(g6758A));
AND2_X1 U_g9713A (.ZN(g9713A),.A2(FE_OFN63_g9474A),.A1(g1589A));
AND2_X1 U_g4431A (.ZN(g4431A),.A2(g3533A),.A1(g2268A));
AND2_X1 U_g4252A (.ZN(g4252A),.A2(FE_OFN347_g3914A),.A1(g1007A));
AND2_X1 U_g11166A (.ZN(g11166A),.A2(FE_OFN9_g10702A),.A1(g542A));
AND2_X1 U_g7130A (.ZN(g7130A),.A2(g6697A),.A1(g5150A));
AND2_X1 U_g11009A (.ZN(g11009A),.A2(FE_OFN18_g10702A),.A1(g5179A));
AND2_X1 U_g7542A (.ZN(g7542A),.A2(g79A),.A1(FE_OFN85_g2176A));
AND2_X1 U_g8019A (.ZN(g8019A),.A2(FE_OFN310_g4336A),.A1(g6573A));
AND2_X1 U_g11008A (.ZN(g11008A),.A2(FE_OFN18_g10702A),.A1(g5171A));
AND2_X1 U_g3516A (.ZN(g3516A),.A2(FE_OFN298_g3015A),.A1(g1209A));
AND2_X1 U_g8052A (.ZN(g8052A),.A2(FE_OFN305_g5151A),.A1(g7573A));
AND2_X1 U_g3987A (.ZN(g3987A),.A2(FE_OFN359_g18A),.A1(g243A));
AND2_X1 U_g4765A (.ZN(g4765A),.A2(FE_OFN307_g4010A),.A1(g491A));
AND2_X1 U_g11555A (.ZN(g11555A),.A2(FE_OFN27_g11519A),.A1(FE_OFN238_g1781A));
AND2_X1 U_g9857A (.ZN(g9857A),.A2(g9569A),.A1(g9734A));
AND2_X1 U_g8728A (.ZN(g8728A),.A2(g7915A),.A1(g8226A));
AND2_X1 U_g8730A (.ZN(g8730A),.A2(g7917A),.A1(g8230A));
AND2_X1 U_g8185A (.ZN(g8185A),.A2(g8234A),.A1(g664A));
AND2_X1 U_g5194A (.ZN(g5194A),.A2(FE_OFN299_g4457A),.A1(g1610A));
AND2_X1 U_g8385A (.ZN(g8385A),.A2(g8234A),.A1(g5255A));
AND2_X1 U_g4610A (.ZN(g4610A),.A2(g2212A),.A1(g3804A));
AND2_X1 U_g7902A (.ZN(g7902A),.A2(g6449A),.A1(g7661A));
AND2_X1 U_g4073A (.ZN(g4073A),.A2(g3222A),.A1(g3200A));
AND2_X1 U_g8070A (.ZN(g8070A),.A2(FE_OFN198_g7697A),.A1(g682A));
AND2_X1 U_g5731A (.ZN(g5731A),.A2(FE_OFN315_g5117A),.A1(g1583A));
AND2_X1 U_g11238A (.ZN(g11238A),.A2(g11111A),.A1(g4553A));
AND2_X1 U_g4473A (.ZN(g4473A),.A2(FE_OFN302_g3913A),.A1(g1125A));
AND2_X1 U_g8470A (.ZN(g8470A),.A2(FE_OFN210_g7246A),.A1(g8308A));
AND2_X1 U_g5489A (.ZN(g5489A),.A2(FE_OFN358_g3521A),.A1(g557A));
AND2_X1 U_g3991A (.ZN(g3991A),.A2(g2774A),.A1(g1738A));
AND4_X1 U_I5887A (.ZN(I5887A),.A4(g2095A),.A3(g166A),.A2(g2083A),.A1(g2078A));
AND2_X1 U_g7823A (.ZN(g7823A),.A2(FE_OFN209_g6863A),.A1(g1923A));
AND2_X1 U_g4069A (.ZN(g4069A),.A2(g2777A),.A1(g1762A));
AND3_X4 U_g11519A (.ZN(g11519A),.A3(g11492A),.A2(g3015A),.A1(g1317A));
AND2_X1 U_g11176A (.ZN(g11176A),.A2(FE_OFN20_g10702A),.A1(g506A));
AND2_X1 U_g11092A (.ZN(g11092A),.A2(FE_OFN4_g10950A),.A1(g837A));
AND2_X1 U_g11154A (.ZN(g11154A),.A2(FE_OFN278_g10927A),.A1(g330A));
AND2_X1 U_g9608A (.ZN(g9608A),.A2(FE_OFN71_g9292A),.A1(g7A));
AND2_X1 U_g11637A (.ZN(g11637A),.A2(FE_OFN99_g4421A),.A1(g11596A));
AND2_X1 U_g2091A (.ZN(g2091A),.A2(g971A),.A1(g976A));
AND2_X1 U_g8406A (.ZN(g8406A),.A2(g8146A),.A1(g695A));
AND2_X1 U_g5254A (.ZN(g5254A),.A2(FE_OFN357_g3521A),.A1(g549A));
AND2_X1 U_g7260A (.ZN(g7260A),.A2(g2345A),.A1(g6752A));
AND2_X1 U_g5150A (.ZN(g5150A),.A2(g4678A),.A1(g1275A));
AND2_X1 U_g8766A (.ZN(g8766A),.A2(FE_OFN304_g5151A),.A1(g8612A));
AND2_X1 U_g9588A (.ZN(g9588A),.A2(FE_OFN53_g9173A),.A1(g1351A));
AND2_X1 U_g8801A (.ZN(g8801A),.A2(FE_OFN331_g8696A),.A1(g8742A));
AND2_X1 U_g7063A (.ZN(g7063A),.A2(g6586A),.A1(g5008A));
AND2_X1 U_g10303A (.ZN(g10303A),.A2(g9291A),.A1(g9995A));
AND2_X1 U_g5009A (.ZN(g5009A),.A2(FE_OFN154_g4640A),.A1(g1486A));
AND2_X1 U_g9665A (.ZN(g9665A),.A2(FE_OFN48_g9151A),.A1(g1314A));
AND2_X2 U_g8748A (.ZN(g8748A),.A2(g8488A),.A1(I9810A));
AND2_X1 U_g11215A (.ZN(g11215A),.A2(FE_OFN279_g11157A),.A1(g953A));
AND2_X1 U_g10750A (.ZN(g10750A),.A2(FE_OFN102_g3586A),.A1(g10597A));
AND3_X1 U_g5769A (.ZN(g5769A),.A3(g3818A),.A2(FE_OFN200_g4921A),.A1(g3092A));
AND2_X1 U_g6673A (.ZN(g6673A),.A2(I9326A),.A1(g90A));
AND2_X1 U_g5212A (.ZN(g5212A),.A2(g4678A),.A1(g1255A));
AND2_X1 U_g7720A (.ZN(g7720A),.A2(FE_OFN191_g6488A),.A1(g727A));
AND3_X1 U_g5918A (.ZN(g5918A),.A3(g4609A),.A2(FE_OFN184_I7048A),.A1(g109A));
AND2_X1 U_g8045A (.ZN(g8045A),.A2(g5128A),.A1(g7547A));
AND2_X1 U_g8173A (.ZN(g8173A),.A2(FE_OFN363_I5565A),.A1(g7971A));
AND2_X1 U_g11349A (.ZN(g11349A),.A2(g7914A),.A1(g11288A));
AND2_X1 U_g7843A (.ZN(g7843A),.A2(g5919A),.A1(g7599A));
AND2_X1 U_g9696A (.ZN(g9696A),.A2(FE_OFN59_g9432A),.A1(g281A));
AND2_X1 U_g6772A (.ZN(g6772A),.A2(g722A),.A1(g6228A));
AND2_X1 U_g6058A (.ZN(g6058A),.A2(g85A),.A1(g1035A));
AND2_X1 U_g6531A (.ZN(g6531A),.A2(FE_OFN283_I8869A),.A1(g79A));
AND2_X1 U_g6743A (.ZN(g6743A),.A2(FE_OFN219_g5557A),.A1(g4106A));
AND2_X1 U_g6890A (.ZN(g6890A),.A2(g6403A),.A1(g6752A));
AND2_X1 U_g7549A (.ZN(g7549A),.A2(FE_OFN137_g3829A),.A1(g7269A));
AND2_X1 U_g8169A (.ZN(g8169A),.A2(I11360A),.A1(g35A));
AND2_X1 U_g11304A (.ZN(g11304A),.A2(g11243A),.A1(g4585A));
AND2_X1 U_g9944A (.ZN(g9944A),.A2(FE_OFN68_g9392A),.A1(g9924A));
AND2_X4 U_g9240A (.ZN(g9240A),.A2(g8962A),.A1(FE_OFN277_g48A));
AND2_X1 U_g8059A (.ZN(g8059A),.A2(FE_OFN177_g5919A),.A1(g7592A));
AND2_X1 U_g8718A (.ZN(g8718A),.A2(g7903A),.A1(g8203A));
AND2_X1 U_g8767A (.ZN(g8767A),.A2(FE_OFN304_g5151A),.A1(g8616A));
AND2_X1 U_g9316A (.ZN(g9316A),.A2(g48A),.A1(g8877A));
AND2_X1 U_g7625A (.ZN(g7625A),.A2(FE_OFN191_g6488A),.A1(g673A));
AND2_X1 U_g8793A (.ZN(g8793A),.A2(FE_OFN331_g8696A),.A1(g8644A));
AND2_X1 U_g2940A (.ZN(g2940A),.A2(g1654A),.A1(g2424A));
AND2_X1 U_g4114A (.ZN(g4114A),.A2(g3301A),.A1(g1351A));
AND2_X1 U_g11636A (.ZN(g11636A),.A2(g7897A),.A1(g11624A));
AND2_X1 U_g10949A (.ZN(g10949A),.A2(g10809A),.A1(g2947A));
AND2_X1 U_g3563A (.ZN(g3563A),.A2(g2126A),.A1(g3275A));
AND2_X1 U_g10948A (.ZN(g10948A),.A2(g10809A),.A1(g2223A));
AND2_X1 U_g8246A (.ZN(g8246A),.A2(g7438A),.A1(g7846A));
AND2_X1 U_g5788A (.ZN(g5788A),.A2(g5222A),.A1(g1540A));
AND2_X1 U_g4008A (.ZN(g4008A),.A2(FE_OFN224_g2276A),.A1(FE_OFN236_g1776A));
AND2_X1 U_g9596A (.ZN(g9596A),.A2(g9010A),.A1(g928A));
AND2_X1 U_g5249A (.ZN(g5249A),.A2(FE_OFN288_g4263A),.A1(g1089A));
AND2_X1 U_g11585A (.ZN(g11585A),.A2(g11539A),.A1(g1321A));
AND2_X1 U_g3089A (.ZN(g3089A),.A2(g2050A),.A1(g2054A));
AND2_X1 U_g4972A (.ZN(g4972A),.A2(FE_OFN147_g4682A),.A1(g1436A));
AND2_X1 U_g11554A (.ZN(g11554A),.A2(FE_OFN27_g11519A),.A1(g1776A));
AND2_X1 U_g7586A (.ZN(g7586A),.A2(g5420A),.A1(g7096A));
AND2_X1 U_g10673A (.ZN(g10673A),.A2(FE_OFN79_g8700A),.A1(g10417A));
AND3_X1 U_g4806A (.ZN(g4806A),.A3(g2493A),.A2(g3992A),.A1(g3215A));
AND2_X1 U_g5485A (.ZN(g5485A),.A2(FE_OFN333_g4294A),.A1(g1914A));
AND2_X1 U_g9936A (.ZN(g9936A),.A2(FE_OFN60_g9624A),.A1(g9915A));
AND2_X1 U_g2910A (.ZN(g2910A),.A2(g1660A),.A1(g2424A));
AND2_X1 U_g9317A (.ZN(g9317A),.A2(g8875A),.A1(g6109A));
AND2_X1 U_g10933A (.ZN(g10933A),.A2(g3982A),.A1(g10853A));
AND2_X1 U_g8388A (.ZN(g8388A),.A2(g7246A),.A1(g8177A));
AND2_X1 U_g4465A (.ZN(g4465A),.A2(FE_OFN302_g3913A),.A1(g1117A));
AND2_X1 U_g7141A (.ZN(g7141A),.A2(g6716A),.A1(g5230A));
AND2_X1 U_g10508A (.ZN(g10508A),.A2(FE_OFN336_g1690A),.A1(g10013A));
AND2_X1 U_g4230A (.ZN(g4230A),.A2(FE_OFN132_g3015A),.A1(g1095A));
AND2_X1 U_g10634A (.ZN(g10634A),.A2(g3829A),.A1(g10382A));
AND2_X1 U_g9601A (.ZN(g9601A),.A2(g9192A),.A1(g922A));
AND2_X1 U_g6126A (.ZN(g6126A),.A2(FE_OFN322_g4449A),.A1(g3681A));
AND2_X1 U_g6326A (.ZN(g6326A),.A2(FE_OFN115_g4807A),.A1(g1250A));
AND2_X1 U_g7710A (.ZN(g7710A),.A2(FE_OFN191_g6488A),.A1(g700A));
AND2_X1 U_g8028A (.ZN(g8028A),.A2(g7438A),.A1(g7375A));
AND2_X1 U_g6760A (.ZN(g6760A),.A2(g6221A),.A1(g786A));
AND2_X1 U_g5640A (.ZN(g5640A),.A2(FE_OFN290_g4880A),.A1(g1059A));
AND2_X1 U_g5031A (.ZN(g5031A),.A2(FE_OFN153_g4640A),.A1(g1478A));
AND2_X1 U_g4550A (.ZN(g4550A),.A2(FE_OFN344_g3586A),.A1(g342A));
AND2_X1 U_g7879A (.ZN(g7879A),.A2(FE_OFN366_g3521A),.A1(g5286A));
AND2_X1 U_g7962A (.ZN(g7962A),.A2(g6403A),.A1(g7730A));
AND2_X1 U_g9597A (.ZN(g9597A),.A2(FE_OFN46_g9125A),.A1(g1170A));
AND2_X1 U_g10452A (.ZN(g10452A),.A2(FE_OFN234_g2024A),.A1(g10439A));
AND2_X1 U_g4891A (.ZN(g4891A),.A2(g4739A),.A1(g631A));
AND2_X1 U_g5005A (.ZN(g5005A),.A2(FE_OFN154_g4640A),.A1(g1490A));
AND2_X1 U_g6423A (.ZN(g6423A),.A2(FE_OFN217_g5013A),.A1(g4348A));
AND2_X1 U_g8108A (.ZN(g8108A),.A2(g7952A),.A1(g1891A));
AND3_X4 U_g4807A (.ZN(g4807A),.A3(I6360A),.A2(g1289A),.A1(g3015A));
AND2_X1 U_g5911A (.ZN(g5911A),.A2(g4977A),.A1(g3322A));
AND2_X1 U_g9937A (.ZN(g9937A),.A2(FE_OFN60_g9624A),.A1(g9916A));
AND2_X1 U_g9840A (.ZN(g9840A),.A2(g9747A),.A1(g9704A));
AND2_X1 U_g10780A (.ZN(g10780A),.A2(g4467A),.A1(g10723A));
AND2_X1 U_g8217A (.ZN(g8217A),.A2(g7883A),.A1(g1872A));
AND2_X1 U_g11013A (.ZN(g11013A),.A2(FE_OFN18_g10702A),.A1(g5209A));
AND2_X1 U_g9390A (.ZN(g9390A),.A2(FE_OFN48_g9151A),.A1(g1333A));
AND2_X1 U_g11214A (.ZN(g11214A),.A2(FE_OFN279_g11157A),.A1(g950A));
AND2_X1 U_g6327A (.ZN(g6327A),.A2(FE_OFN115_g4807A),.A1(g1255A));
AND2_X1 U_g4342A (.ZN(g4342A),.A2(FE_OFN351_g3913A),.A1(g1149A));
AND2_X1 U_g5796A (.ZN(g5796A),.A2(FE_OFN321_g5261A),.A1(g1564A));
AND2_X1 U_g5473A (.ZN(g5473A),.A2(FE_OFN367_g3521A),.A1(g546A));
AND2_X1 U_g6346A (.ZN(g6346A),.A2(g5878A),.A1(g5038A));
AND2_X1 U_g6633A (.ZN(g6633A),.A2(FE_OFN282_g6165A),.A1(g354A));
AND2_X1 U_g11005A (.ZN(g11005A),.A2(FE_OFN13_g10702A),.A1(g5119A));
AND2_X1 U_g8365A (.ZN(g8365A),.A2(g8146A),.A1(g668A));
AND2_X1 U_g8048A (.ZN(g8048A),.A2(g5919A),.A1(g7558A));
AND2_X1 U_g4481A (.ZN(g4481A),.A2(g3906A),.A1(g1713A));
AND2_X1 U_g4097A (.ZN(g4097A),.A2(g3060A),.A1(g2677A));
AND2_X1 U_g8055A (.ZN(g8055A),.A2(FE_OFN305_g5151A),.A1(g7588A));
AND2_X1 U_g4497A (.ZN(g4497A),.A2(FE_OFN344_g3586A),.A1(g351A));
AND2_X1 U_g9942A (.ZN(g9942A),.A2(FE_OFN67_g9367A),.A1(g9922A));
AND2_X1 U_g6696A (.ZN(g6696A),.A2(I9326A),.A1(g94A));
AND3_X1 U_g10731A (.ZN(g10731A),.A3(g10665A),.A2(g1850A),.A1(g5118A));
AND2_X1 U_g8827A (.ZN(g8827A),.A2(g8696A),.A1(g8552A));
AND2_X1 U_g5540A (.ZN(g5540A),.A2(g4292A),.A1(g1727A));
AND2_X1 U_g4960A (.ZN(g4960A),.A2(FE_OFN147_g4682A),.A1(g1403A));
AND2_X1 U_g8846A (.ZN(g8846A),.A2(FE_OFN328_g8709A),.A1(g8615A));
AND2_X1 U_g6508A (.ZN(g6508A),.A2(FE_OFN363_I5565A),.A1(g5983A));
AND2_X1 U_g6240A (.ZN(g6240A),.A2(g5361A),.A1(g182A));
AND2_X1 U_g7931A (.ZN(g7931A),.A2(g7446A),.A1(g52A));
AND2_X1 U_g5287A (.ZN(g5287A),.A2(g4782A),.A1(I6260A));
AND2_X1 U_g6472A (.ZN(g6472A),.A2(g1936A),.A1(g5853A));
AND2_X1 U_g11100A (.ZN(g11100A),.A2(FE_OFN4_g10950A),.A1(g853A));
AND2_X1 U_g11235A (.ZN(g11235A),.A2(g11107A),.A1(g4529A));
AND2_X1 U_g5199A (.ZN(g5199A),.A2(FE_OFN288_g4263A),.A1(g1068A));
AND2_X1 U_g6316A (.ZN(g6316A),.A2(FE_OFN117_g4807A),.A1(g1270A));
AND2_X1 U_g7515A (.ZN(g7515A),.A2(g70A),.A1(FE_OFN85_g2176A));
AND2_X1 U_g10583A (.ZN(g10583A),.A2(g10515A),.A1(g10518A));
AND2_X1 U_g5781A (.ZN(g5781A),.A2(g5222A),.A1(g1537A));
AND2_X1 U_g8018A (.ZN(g8018A),.A2(g7438A),.A1(g7742A));
AND2_X1 U_g4401A (.ZN(g4401A),.A2(g3772A),.A1(g1845A));
AND3_X1 U_g8994A (.ZN(g8994A),.A3(g8783A),.A2(FE_OFN92_g2216A),.A1(g8110A));
AND2_X1 U_g2950A (.ZN(g2950A),.A2(g1666A),.A1(g2424A));
AND2_X1 U_g5510A (.ZN(g5510A),.A2(g4289A),.A1(g1630A));
AND2_X1 U_g6347A (.ZN(g6347A),.A2(FE_OFN320_g5361A),.A1(g275A));
AND2_X1 U_g9357A (.ZN(g9357A),.A2(g9223A),.A1(g962A));
AND2_X1 U_g4828A (.ZN(g4828A),.A2(g695A),.A1(g4106A));
AND2_X1 U_g11407A (.ZN(g11407A),.A2(g4807A),.A1(g11249A));
AND2_X1 U_g4727A (.ZN(g4727A),.A2(FE_OFN300_g4002A),.A1(g386A));
AND2_X1 U_g10357A (.ZN(g10357A),.A2(FE_OFN269_g109A),.A1(I15500A));
AND2_X1 U_g10743A (.ZN(g10743A),.A2(FE_OFN364_g3015A),.A1(g10639A));
AND2_X1 U_g5259A (.ZN(g5259A),.A2(g4739A),.A1(g627A));
AND2_X1 U_g5694A (.ZN(g5694A),.A2(FE_OFN365_g5361A),.A1(g162A));
AND2_X1 U_g10769A (.ZN(g10769A),.A2(FE_OFN297_g3015A),.A1(g10652A));
AND2_X1 U_g11584A (.ZN(g11584A),.A2(g11539A),.A1(g1318A));
AND2_X1 U_g4932A (.ZN(g4932A),.A2(FE_OFN290_g4880A),.A1(g1065A));
AND2_X1 U_g10768A (.ZN(g10768A),.A2(FE_OFN293_g3015A),.A1(g10649A));
AND2_X1 U_g6820A (.ZN(g6820A),.A2(FE_OFN178_g5354A),.A1(g1362A));
AND2_X1 U_g4068A (.ZN(g4068A),.A2(FE_OFN224_g2276A),.A1(FE_OFN251_g1801A));
AND2_X1 U_g6317A (.ZN(g6317A),.A2(FE_OFN117_g4807A),.A1(g1304A));
AND2_X1 U_g5215A (.ZN(g5215A),.A2(g3275A),.A1(g4276A));
AND2_X1 U_g4576A (.ZN(g4576A),.A2(g4010A),.A1(g530A));
AND2_X1 U_g6775A (.ZN(g6775A),.A2(g6231A),.A1(g822A));
AND2_X4 U_g3829A (.ZN(g3829A),.A2(g1696A),.A1(g2028A));
AND2_X1 U_g10662A (.ZN(g10662A),.A2(g10396A),.A1(g8700A));
AND2_X1 U_g8101A (.ZN(g8101A),.A2(FE_OFN207_g6863A),.A1(g5484A));
AND2_X1 U_g5825A (.ZN(g5825A),.A2(g5318A),.A1(g3204A));
AND4_X1 U_I6310A (.ZN(I6310A),.A4(g2435A),.A3(g2421A),.A2(g2407A),.A1(g2396A));
AND2_X1 U_g7884A (.ZN(g7884A),.A2(FE_OFN334_g7045A),.A1(g7457A));
AND2_X1 U_g5008A (.ZN(g5008A),.A2(FE_OFN303_g4678A),.A1(g1292A));
AND2_X1 U_g3974A (.ZN(g3974A),.A2(FE_OFN260_g18A),.A1(g231A));
AND2_X1 U_g9949A (.ZN(g9949A),.A2(FE_OFN68_g9392A),.A1(g9929A));
AND2_X1 U_g2531A (.ZN(g2531A),.A2(g668A),.A1(g658A));
AND2_X2 U_g9292A (.ZN(g9292A),.A2(g48A),.A1(g8878A));
AND2_X1 U_g10778A (.ZN(g10778A),.A2(g10679A),.A1(g1027A));
AND2_X1 U_g8041A (.ZN(g8041A),.A2(g5128A),.A1(g7524A));
AND2_X1 U_g6079A (.ZN(g6079A),.A2(FE_OFN273_g85A),.A1(g1053A));
AND2_X1 U_g7235A (.ZN(g7235A),.A2(g6447A),.A1(g6663A));
AND2_X1 U_g9603A (.ZN(g9603A),.A2(FE_OFN46_g9125A),.A1(g1173A));
AND2_X1 U_g6840A (.ZN(g6840A),.A2(FE_OFN180_g5354A),.A1(g248A));
AND2_X1 U_g9850A (.ZN(g9850A),.A2(g9579A),.A1(g9726A));
AND2_X1 U_g7988A (.ZN(g7988A),.A2(g7379A),.A1(g1878A));
AND2_X1 U_g5228A (.ZN(g5228A),.A2(FE_OFN288_g4263A),.A1(g1086A));
AND2_X1 U_g7134A (.ZN(g7134A),.A2(g6354A),.A1(g5587A));
AND2_X1 U_g5934A (.ZN(g5934A),.A2(g1965A),.A1(g5215A));
AND2_X1 U_g5230A (.ZN(g5230A),.A2(g4678A),.A1(g1265A));
AND2_X1 U_g8168A (.ZN(g8168A),.A2(FE_OFN89_I11360A),.A1(g34A));
AND2_X1 U_g9583A (.ZN(g9583A),.A2(g8995A),.A1(g886A));
AND2_X1 U_g10672A (.ZN(g10672A),.A2(g9473A),.A1(g10414A));
AND2_X1 U_g3287A (.ZN(g3287A),.A2(g5188A),.A1(g802A));
AND2_X1 U_g8772A (.ZN(g8772A),.A2(FE_OFN304_g5151A),.A1(g8627A));
AND2_X1 U_g4893A (.ZN(g4893A),.A2(g4739A),.A1(g635A));
AND2_X1 U_g10331A (.ZN(g10331A),.A2(FE_OFN269_g109A),.A1(I15510A));
AND2_X1 U_g8505A (.ZN(g8505A),.A2(FE_OFN359_g18A),.A1(g8309A));
AND2_X1 U_g10449A (.ZN(g10449A),.A2(FE_OFN235_g2024A),.A1(g10433A));
AND2_X1 U_g11273A (.ZN(g11273A),.A2(g11199A),.A1(g4765A));
AND2_X1 U_g8734A (.ZN(g8734A),.A2(g7923A),.A1(g8187A));
AND2_X1 U_g5913A (.ZN(g5913A),.A2(g85A),.A1(g1041A));
AND2_X1 U_g10448A (.ZN(g10448A),.A2(FE_OFN235_g2024A),.A1(g10421A));
AND2_X1 U_g6163A (.ZN(g6163A),.A2(g5354A),.A1(g4572A));
AND2_X1 U_g6363A (.ZN(g6363A),.A2(FE_OFN320_g5361A),.A1(g284A));
AND2_X1 U_g7202A (.ZN(g7202A),.A2(FE_OFN322_g4449A),.A1(g5226A));
AND2_X1 U_g11463A (.ZN(g11463A),.A2(FE_OFN99_g4421A),.A1(g11229A));
AND2_X1 U_g8074A (.ZN(g8074A),.A2(FE_OFN198_g7697A),.A1(g718A));
AND2_X1 U_g4325A (.ZN(g4325A),.A2(FE_OFN351_g3913A),.A1(g1166A));
AND2_X1 U_g8474A (.ZN(g8474A),.A2(g5521A),.A1(g8383A));
AND2_X1 U_g11234A (.ZN(g11234A),.A2(g11107A),.A1(g4518A));
AND2_X1 U_g5266A (.ZN(g5266A),.A2(FE_OFN335_g4737A),.A1(g718A));
AND2_X1 U_g4483A (.ZN(g4483A),.A2(FE_OFN103_g3586A),.A1(g336A));
AND2_X1 U_g5248A (.ZN(g5248A),.A2(FE_OFN335_g4737A),.A1(g673A));
AND2_X1 U_g11514A (.ZN(g11514A),.A2(FE_OFN176_g5151A),.A1(g11491A));
AND2_X1 U_g5255A (.ZN(g5255A),.A2(FE_OFN335_g4737A),.A1(g682A));
AND2_X1 U_g4106A (.ZN(g4106A),.A2(g686A),.A1(g3284A));
AND2_X1 U_g2760A (.ZN(g2760A),.A2(g2091A),.A1(g981A));
AND2_X1 U_g5097A (.ZN(g5097A),.A2(g4608A),.A1(g1786A));
AND2_X1 U_g5726A (.ZN(g5726A),.A2(FE_OFN315_g5117A),.A1(g1601A));
AND2_X1 U_g5497A (.ZN(g5497A),.A2(FE_OFN357_g3521A),.A1(g560A));
AND2_X4 U_g5354A (.ZN(g5354A),.A2(I7048A),.A1(FE_OFN352_g109A));
AND2_X1 U_g7933A (.ZN(g7933A),.A2(g7450A),.A1(g55A));
AND2_X1 U_g9617A (.ZN(g9617A),.A2(g9274A),.A1(g9A));
AND2_X1 U_g9906A (.ZN(g9906A),.A2(g9680A),.A1(g9873A));
AND2_X1 U_g11012A (.ZN(g11012A),.A2(FE_OFN18_g10702A),.A1(g5196A));
AND2_X1 U_g7050A (.ZN(g7050A),.A2(g6702A),.A1(g5001A));
AND2_X1 U_g10971A (.ZN(g10971A),.A2(g2045A),.A1(g10849A));
AND2_X1 U_g4904A (.ZN(g4904A),.A2(g4243A),.A1(g1850A));
AND2_X1 U_g10369A (.ZN(g10369A),.A2(FE_OFN235_g2024A),.A1(g10361A));
AND2_X1 U_g8400A (.ZN(g8400A),.A2(g8234A),.A1(g5271A));
AND2_X1 U_g4345A (.ZN(g4345A),.A2(FE_OFN289_g4679A),.A1(g1169A));
AND2_X1 U_g2161A (.ZN(g2161A),.A2(I5085A),.A1(I5084A));
AND2_X1 U_g5001A (.ZN(g5001A),.A2(FE_OFN303_g4678A),.A1(g1300A));
AND2_X1 U_g9945A (.ZN(g9945A),.A2(FE_OFN68_g9392A),.A1(g9925A));
AND2_X1 U_g7271A (.ZN(g7271A),.A2(g6354A),.A1(g5028A));
AND2_X1 U_g9709A (.ZN(g9709A),.A2(FE_OFN70_g9490A),.A1(g1524A));
AND2_X1 U_g4223A (.ZN(g4223A),.A2(FE_OFN347_g3914A),.A1(g1003A));
AND2_X1 U_g10716A (.ZN(g10716A),.A2(g10396A),.A1(g10497A));
AND2_X1 U_g11291A (.ZN(g11291A),.A2(g4379A),.A1(g11247A));
AND2_X1 U_g6661A (.ZN(g6661A),.A2(FE_OFN97_I8869A),.A1(g73A));
AND2_X1 U_g11173A (.ZN(g11173A),.A2(FE_OFN21_g10702A),.A1(g491A));
AND2_X1 U_g6075A (.ZN(g6075A),.A2(g5613A),.A1(g549A));
AND2_X1 U_g8023A (.ZN(g8023A),.A2(g7438A),.A1(g7367A));
AND2_X1 U_g9907A (.ZN(g9907A),.A2(g9680A),.A1(g9888A));
AND2_X1 U_g10582A (.ZN(g10582A),.A2(g9473A),.A1(g10339A));
AND2_X1 U_g5746A (.ZN(g5746A),.A2(FE_OFN353_g5117A),.A1(g1589A));
AND2_X1 U_g5221A (.ZN(g5221A),.A2(g4678A),.A1(g1260A));
AND2_X1 U_g9959A (.ZN(g9959A),.A2(FE_OFN280_g9536A),.A1(g9950A));
AND2_X1 U_g7674A (.ZN(g7674A),.A2(g3880A),.A1(g5857A));
AND2_X1 U_g9690A (.ZN(g9690A),.A2(g9432A),.A1(g266A));
AND2_X1 U_g6627A (.ZN(g6627A),.A2(FE_OFN283_I8869A),.A1(g58A));
AND2_X1 U_g5703A (.ZN(g5703A),.A2(FE_OFN365_g5361A),.A1(g174A));
AND2_X1 U_g4522A (.ZN(g4522A),.A2(FE_OFN344_g3586A),.A1(g360A));
AND2_X1 U_g4115A (.ZN(g4115A),.A2(g3060A),.A1(FE_OFN236_g1776A));
AND2_X1 U_g7541A (.ZN(g7541A),.A2(I6360A),.A1(g7075A));
AND2_X1 U_g10627A (.ZN(g10627A),.A2(FE_OFN227_g3880A),.A1(g10452A));
AND2_X1 U_g4047A (.ZN(g4047A),.A2(FE_OFN225_g2276A),.A1(FE_OFN238_g1781A));
AND2_X1 U_g6526A (.ZN(g6526A),.A2(FE_OFN283_I8869A),.A1(g76A));
AND2_X1 U_g2944A (.ZN(g2944A),.A2(g1669A),.A1(g2424A));
AND2_X1 U_g6646A (.ZN(g6646A),.A2(g6165A),.A1(g360A));
AND2_X1 U_g7132A (.ZN(g7132A),.A2(g6702A),.A1(g5182A));
AND2_X1 U_g11029A (.ZN(g11029A),.A2(FE_OFN17_g10702A),.A1(g401A));
AND2_X1 U_g8051A (.ZN(g8051A),.A2(FE_OFN305_g5151A),.A1(g7572A));
AND2_X1 U_g8127A (.ZN(g8127A),.A2(g7949A),.A1(g1927A));
AND2_X1 U_g7209A (.ZN(g7209A),.A2(g6432A),.A1(g3804A));
AND2_X1 U_g11028A (.ZN(g11028A),.A2(FE_OFN17_g10702A),.A1(g396A));
AND2_X1 U_g6439A (.ZN(g6439A),.A2(g5919A),.A1(g3631A));
AND2_X1 U_g10742A (.ZN(g10742A),.A2(g3586A),.A1(g10655A));
AND2_X1 U_g9110A (.ZN(g9110A),.A2(FE_OFN359_g18A),.A1(g8880A));
AND2_X1 U_g10681A (.ZN(g10681A),.A2(g3586A),.A1(g10567A));
AND2_X1 U_g4537A (.ZN(g4537A),.A2(g4002A),.A1(g444A));
AND2_X1 U_g9663A (.ZN(g9663A),.A2(FE_OFN39_g9223A),.A1(g959A));
AND2_X1 U_g5349A (.ZN(g5349A),.A2(g4617A),.A1(g2126A));
AND2_X1 U_g8732A (.ZN(g8732A),.A2(g7919A),.A1(g8200A));
AND2_X1 U_g3807A (.ZN(g3807A),.A2(g3062A),.A1(g3003A));
AND2_X1 U_g5848A (.ZN(g5848A),.A2(g5519A),.A1(g3860A));
AND2_X1 U_g8508A (.ZN(g8508A),.A2(FE_OFN330_g7638A),.A1(g8411A));
AND2_X1 U_g8072A (.ZN(g8072A),.A2(FE_OFN199_g7697A),.A1(g700A));
AND2_X1 U_g5699A (.ZN(g5699A),.A2(g5117A),.A1(g1592A));
AND2_X1 U_g11240A (.ZN(g11240A),.A2(g11111A),.A1(g4560A));
AND2_X1 U_g5398A (.ZN(g5398A),.A2(g2224A),.A1(g4610A));
AND2_X1 U_g6616A (.ZN(g6616A),.A2(FE_OFN363_I5565A),.A1(g6105A));
AND2_X1 U_g10690A (.ZN(g10690A),.A2(FE_OFN136_g3863A),.A1(g10387A));
AND2_X1 U_g8043A (.ZN(g8043A),.A2(FE_OFN305_g5151A),.A1(g7582A));
AND2_X1 U_g9590A (.ZN(g9590A),.A2(g8995A),.A1(g895A));
AND2_X1 U_g4128A (.ZN(g4128A),.A2(g627A),.A1(g1976A));
AND2_X1 U_g6404A (.ZN(g6404A),.A2(FE_OFN217_g5013A),.A1(g2132A));
AND2_X1 U_g6647A (.ZN(g6647A),.A2(g5808A),.A1(g87A));
AND2_X1 U_g10504A (.ZN(g10504A),.A2(FE_OFN336_g1690A),.A1(g10001A));
AND2_X1 U_g9657A (.ZN(g9657A),.A2(g9205A),.A1(g919A));
AND2_X1 U_g4542A (.ZN(g4542A),.A2(FE_OFN344_g3586A),.A1(g366A));
AND2_X1 U_g4330A (.ZN(g4330A),.A2(FE_OFN351_g3913A),.A1(g1163A));
AND2_X1 U_g3497A (.ZN(g3497A),.A2(g1900A),.A1(g2804A));
AND2_X1 U_g5524A (.ZN(g5524A),.A2(g3906A),.A1(g1678A));
AND2_X1 U_g8147A (.ZN(g8147A),.A2(g7907A),.A1(g928A));
AND2_X1 U_g4554A (.ZN(g4554A),.A2(g4010A),.A1(g542A));
AND2_X1 U_g9899A (.ZN(g9899A),.A2(g9367A),.A1(g9713A));
AND2_X1 U_g5258A (.ZN(g5258A),.A2(FE_OFN335_g4737A),.A1(g700A));
AND2_X1 U_g7736A (.ZN(g7736A),.A2(FE_OFN226_g3880A),.A1(g5814A));
AND2_X1 U_g6224A (.ZN(g6224A),.A2(FE_OFN306_g5128A),.A1(g1520A));
AND2_X1 U_g10626A (.ZN(g10626A),.A2(FE_OFN369_g4525A),.A1(g10453A));
AND2_X1 U_g6320A (.ZN(g6320A),.A2(FE_OFN118_g4807A),.A1(g1292A));
AND2_X1 U_g7623A (.ZN(g7623A),.A2(FE_OFN191_g6488A),.A1(g664A));
AND2_X1 U_g10299A (.ZN(g10299A),.A2(g10013A),.A1(FE_OFN76_g8700A));
AND2_X1 U_g7889A (.ZN(g7889A),.A2(g3814A),.A1(g5304A));
AND2_X1 U_g10298A (.ZN(g10298A),.A2(g10007A),.A1(g8700A));
AND2_X1 U_g8413A (.ZN(g8413A),.A2(g8146A),.A1(g722A));
AND2_X1 U_g3979A (.ZN(g3979A),.A2(FE_OFN260_g18A),.A1(g237A));
AND2_X1 U_g4902A (.ZN(g4902A),.A2(g4243A),.A1(g1848A));
AND2_X1 U_g5211A (.ZN(g5211A),.A2(FE_OFN288_g4263A),.A1(g1080A));
AND2_X1 U_g4512A (.ZN(g4512A),.A2(FE_OFN344_g3586A),.A1(g357A));
AND2_X1 U_g7722A (.ZN(g7722A),.A2(g6449A),.A1(g7127A));
AND2_X1 U_g9844A (.ZN(g9844A),.A2(g9522A),.A1(g9714A));
AND2_X1 U_g4490A (.ZN(g4490A),.A2(FE_OFN302_g3913A),.A1(g1141A));
AND2_X1 U_g6516A (.ZN(g6516A),.A2(FE_OFN363_I5565A),.A1(g5993A));
AND2_X1 U_g5026A (.ZN(g5026A),.A2(FE_OFN153_g4640A),.A1(g1453A));
AND2_X1 U_g8820A (.ZN(g8820A),.A2(g4737A),.A1(g8705A));
AND2_X1 U_g10737A (.ZN(g10737A),.A2(FE_OFN133_g3015A),.A1(g10597A));
AND3_X1 U_g8936A (.ZN(g8936A),.A3(g8849A),.A2(FE_OFN93_g2216A),.A1(g8115A));
AND2_X1 U_g10232A (.ZN(g10232A),.A2(g9974A),.A1(FE_OFN76_g8700A));
AND2_X1 U_g6771A (.ZN(g6771A),.A2(FE_OFN320_g5361A),.A1(g263A));
AND2_X1 U_g5170A (.ZN(g5170A),.A2(g4457A),.A1(g1811A));
AND2_X1 U_g8117A (.ZN(g8117A),.A2(FE_OFN207_g6863A),.A1(g5514A));
AND2_X1 U_g4529A (.ZN(g4529A),.A2(g4002A),.A1(g448A));
AND2_X1 U_g4348A (.ZN(g4348A),.A2(g1909A),.A1(g3497A));
AND2_X1 U_g9966A (.ZN(g9966A),.A2(FE_OFN280_g9536A),.A1(g9956A));
AND2_X1 U_g5280A (.ZN(g5280A),.A2(g2118A),.A1(g3967A));
AND2_X1 U_g7139A (.ZN(g7139A),.A2(g6716A),.A1(g5212A));
AND2_X1 U_g11099A (.ZN(g11099A),.A2(g10883A),.A1(g382A));
AND2_X1 U_g6892A (.ZN(g6892A),.A2(g5013A),.A1(g6472A));
AND2_X1 U_g9705A (.ZN(g9705A),.A2(g9474A),.A1(g1580A));
AND2_X1 U_g10512A (.ZN(g10512A),.A2(FE_OFN336_g1690A),.A1(g10025A));
AND2_X1 U_g11098A (.ZN(g11098A),.A2(FE_OFN4_g10950A),.A1(g849A));
AND2_X1 U_g8775A (.ZN(g8775A),.A2(FE_OFN304_g5151A),.A1(g8628A));
AND2_X1 U_g5083A (.ZN(g5083A),.A2(g4782A),.A1(g2510A));
AND2_X1 U_g5544A (.ZN(g5544A),.A2(FE_OFN291_g4880A),.A1(g1687A));
AND2_X1 U_g11272A (.ZN(g11272A),.A2(g11199A),.A1(g4760A));
AND2_X1 U_g5483A (.ZN(g5483A),.A2(g3906A),.A1(g1621A));
AND2_X1 U_g9948A (.ZN(g9948A),.A2(FE_OFN68_g9392A),.A1(g9928A));
AND2_X1 U_g4063A (.ZN(g4063A),.A2(FE_OFN224_g2276A),.A1(FE_OFN239_g1796A));
AND2_X1 U_g11462A (.ZN(g11462A),.A2(FE_OFN99_g4421A),.A1(g11227A));
AND2_X1 U_g6738A (.ZN(g6738A),.A2(FE_OFN219_g5557A),.A1(g2531A));
AND2_X1 U_g8060A (.ZN(g8060A),.A2(FE_OFN177_g5919A),.A1(g7593A));
AND2_X1 U_g6244A (.ZN(g6244A),.A2(FE_OFN306_g5128A),.A1(g1411A));
AND2_X1 U_g11032A (.ZN(g11032A),.A2(FE_OFN14_g10702A),.A1(g416A));
AND2_X1 U_g10445A (.ZN(g10445A),.A2(g1690A),.A1(g9974A));
AND2_X1 U_g9150A (.ZN(g9150A),.A2(FE_OFN325_g18A),.A1(g8882A));
AND2_X1 U_g10316A (.ZN(g10316A),.A2(g9097A),.A1(g10025A));
AND2_X1 U_g5756A (.ZN(g5756A),.A2(g5261A),.A1(g1531A));
AND2_X1 U_g4720A (.ZN(g4720A),.A2(g4673A),.A1(g1023A));
AND2_X1 U_g9409A (.ZN(g9409A),.A2(g9052A),.A1(g1721A));
AND2_X4 U_g8995A (.ZN(g8995A),.A2(g8929A),.A1(FE_OFN277_g48A));
AND2_X1 U_g6876A (.ZN(g6876A),.A2(g6557A),.A1(g4070A));
AND2_X1 U_g4989A (.ZN(g4989A),.A2(FE_OFN146_g4682A),.A1(g1424A));
AND2_X1 U_g9836A (.ZN(g9836A),.A2(FE_OFN34_g9785A),.A1(g9737A));
AND3_X1 U_g6656A (.ZN(g6656A),.A3(FE_OFN184_I7048A),.A2(g6061A),.A1(g109A));
AND2_X1 U_g5514A (.ZN(g5514A),.A2(FE_OFN333_g4294A),.A1(g1941A));
AND2_X1 U_g8390A (.ZN(g8390A),.A2(g6465A),.A1(g8268A));
AND2_X1 U_g5003A (.ZN(g5003A),.A2(FE_OFN154_g4640A),.A1(g1466A));
AND2_X1 U_g9967A (.ZN(g9967A),.A2(FE_OFN280_g9536A),.A1(g9957A));
AND2_X1 U_g5145A (.ZN(g5145A),.A2(g4673A),.A1(g1639A));
AND2_X1 U_g4971A (.ZN(g4971A),.A2(FE_OFN146_g4682A),.A1(g1419A));
AND2_X1 U_g10753A (.ZN(g10753A),.A2(FE_OFN133_g3015A),.A1(g10649A));
AND2_X1 U_g5695A (.ZN(g5695A),.A2(FE_OFN356_g5361A),.A1(g166A));
AND2_X1 U_g7613A (.ZN(g7613A),.A2(g5013A),.A1(g6940A));
AND2_X1 U_g10736A (.ZN(g10736A),.A2(FE_OFN293_g3015A),.A1(g10658A));
AND2_X1 U_g11220A (.ZN(g11220A),.A2(FE_OFN279_g11157A),.A1(g962A));
AND2_X1 U_g7444A (.ZN(g7444A),.A2(g5557A),.A1(g7277A));
AND2_X1 U_g5536A (.ZN(g5536A),.A2(FE_OFN310_g4336A),.A1(g2970A));
AND2_X1 U_g6663A (.ZN(g6663A),.A2(g2237A),.A1(g6064A));
AND2_X1 U_g4670A (.ZN(g4670A),.A2(g2355A),.A1(g192A));
AND2_X1 U_g6824A (.ZN(g6824A),.A2(FE_OFN178_g5354A),.A1(g1371A));
AND2_X1 U_g4253A (.ZN(g4253A),.A2(FE_OFN132_g3015A),.A1(g1074A));
AND2_X1 U_g8250A (.ZN(g8250A),.A2(g7907A),.A1(g932A));
AND2_X1 U_g8163A (.ZN(g8163A),.A2(g3737A),.A1(g7960A));
AND2_X1 U_g10764A (.ZN(g10764A),.A2(FE_OFN345_g3015A),.A1(g10643A));
AND2_X1 U_g5757A (.ZN(g5757A),.A2(g5222A),.A1(g1552A));
AND2_X1 U_g8032A (.ZN(g8032A),.A2(g7438A),.A1(g7385A));
AND2_X1 U_g11591A (.ZN(g11591A),.A2(g11561A),.A1(g2988A));
AND2_X1 U_g8053A (.ZN(g8053A),.A2(FE_OFN177_g5919A),.A1(g7583A));
AND2_X1 U_g11147A (.ZN(g11147A),.A2(FE_OFN278_g10927A),.A1(g321A));
AND2_X1 U_g5522A (.ZN(g5522A),.A2(g4289A),.A1(g1633A));
AND2_X1 U_g5115A (.ZN(g5115A),.A2(g4572A),.A1(g1394A));
AND2_X1 U_g9837A (.ZN(g9837A),.A2(g9751A),.A1(g9697A));
AND2_X1 U_g9620A (.ZN(g9620A),.A2(FE_OFN40_g9240A),.A1(g976A));
AND2_X1 U_g11151A (.ZN(g11151A),.A2(FE_OFN278_g10927A),.A1(g327A));
AND2_X1 U_g11172A (.ZN(g11172A),.A2(FE_OFN21_g10702A),.A1(g486A));
AND2_X1 U_g7885A (.ZN(g7885A),.A2(g3814A),.A1(g5300A));
AND2_X1 U_g6064A (.ZN(g6064A),.A2(g2230A),.A1(g5398A));
AND3_X1 U_g8929A (.ZN(g8929A),.A3(g8828A),.A2(FE_OFN95_g2216A),.A1(g8095A));
AND2_X1 U_g5595A (.ZN(g5595A),.A2(FE_OFN367_g3521A),.A1(g1621A));
AND2_X1 U_g5537A (.ZN(g5537A),.A2(g4449A),.A1(g2260A));
AND2_X1 U_g9842A (.ZN(g9842A),.A2(g9516A),.A1(g9708A));
AND2_X1 U_g4141A (.ZN(g4141A),.A2(g3060A),.A1(FE_OFN252_g1791A));
AND2_X1 U_g4341A (.ZN(g4341A),.A2(FE_OFN103_g3586A),.A1(g339A));
AND2_X4 U_g9192A (.ZN(g9192A),.A2(g8955A),.A1(FE_OFN277_g48A));
AND2_X1 U_g7679A (.ZN(g7679A),.A2(g6863A),.A1(g1950A));
AND2_X1 U_g7378A (.ZN(g7378A),.A2(FE_OFN226_g3880A),.A1(g5847A));
AND2_X1 U_g5612A (.ZN(g5612A),.A2(FE_OFN357_g3521A),.A1(g1627A));
AND2_X1 U_g7135A (.ZN(g7135A),.A2(g6355A),.A1(g869A));
AND2_X1 U_g10970A (.ZN(g10970A),.A2(g3390A),.A1(g10852A));
AND2_X1 U_g11025A (.ZN(g11025A),.A2(FE_OFN9_g10702A),.A1(g426A));
AND2_X1 U_g9854A (.ZN(g9854A),.A2(g9563A),.A1(g9730A));
AND2_X1 U_g7182A (.ZN(g7182A),.A2(FE_OFN213_g6003A),.A1(g1878A));
AND2_X1 U_g9941A (.ZN(g9941A),.A2(FE_OFN67_g9367A),.A1(g9921A));
AND2_X1 U_g6194A (.ZN(g6194A),.A2(FE_OFN289_g4679A),.A1(g554A));
AND2_X2 U_g5128A (.ZN(g5128A),.A2(FE_OFN352_g109A),.A1(I7048A));
AND2_X1 U_g4962A (.ZN(g4962A),.A2(g4467A),.A1(g1651A));
AND2_X1 U_g4358A (.ZN(g4358A),.A2(g3906A),.A1(g1209A));
AND2_X1 U_g8683A (.ZN(g8683A),.A2(g8549A),.A1(g4803A));
AND2_X1 U_g4506A (.ZN(g4506A),.A2(FE_OFN351_g3913A),.A1(g1113A));
AND2_X1 U_g6471A (.ZN(g6471A),.A2(g5878A),.A1(g5224A));
AND2_X1 U_g8778A (.ZN(g8778A),.A2(g1975A),.A1(g8688A));
AND2_X1 U_g11281A (.ZN(g11281A),.A2(g11203A),.A1(g4788A));
AND2_X1 U_g11146A (.ZN(g11146A),.A2(FE_OFN278_g10927A),.A1(g318A));
AND2_X1 U_g3904A (.ZN(g3904A),.A2(g627A),.A1(g2948A));
AND2_X1 U_g8075A (.ZN(g8075A),.A2(g7697A),.A1(g727A));
AND2_X1 U_g9829A (.ZN(g9829A),.A2(FE_OFN34_g9785A),.A1(g9723A));
AND3_X1 U_g8949A (.ZN(g8949A),.A3(g8828A),.A2(FE_OFN92_g2216A),.A1(g8255A));
AND2_X1 U_g7632A (.ZN(g7632A),.A2(g5420A),.A1(g7184A));
AND2_X1 U_g11290A (.ZN(g11290A),.A2(g4379A),.A1(g11246A));
AND2_X1 U_g6350A (.ZN(g6350A),.A2(FE_OFN346_g4381A),.A1(g5837A));
AND2_X1 U_g10599A (.ZN(g10599A),.A2(g4365A),.A1(g10448A));
AND2_X1 U_g5902A (.ZN(g5902A),.A2(g4977A),.A1(g2555A));
AND4_X1 U_I6337A (.ZN(I6337A),.A4(g2396A),.A3(g2407A),.A2(g2421A),.A1(g201A));
AND2_X2 U_g2276A (.ZN(g2276A),.A2(g1610A),.A1(g1765A));
AND2_X1 U_g6438A (.ZN(g6438A),.A2(g5013A),.A1(g5853A));
AND2_X1 U_g5512A (.ZN(g5512A),.A2(g4281A),.A1(g1660A));
AND2_X1 U_g5090A (.ZN(g5090A),.A2(FE_OFN299_g4457A),.A1(g1781A));
AND2_X1 U_g7719A (.ZN(g7719A),.A2(FE_OFN191_g6488A),.A1(g718A));
AND2_X1 U_g2561A (.ZN(g2561A),.A2(g741A),.A1(g742A));
AND2_X1 U_g3695A (.ZN(g3695A),.A2(FE_OFN292_g3015A),.A1(g1712A));
AND2_X1 U_g8603A (.ZN(g8603A),.A2(g8548A),.A1(g3983A));
AND2_X1 U_g8039A (.ZN(g8039A),.A2(FE_OFN305_g5151A),.A1(g7587A));
AND2_X1 U_g9610A (.ZN(g9610A),.A2(g9192A),.A1(g925A));
AND2_X1 U_g3536A (.ZN(g3536A),.A2(g3103A),.A1(g1289A));
AND2_X1 U_g5529A (.ZN(g5529A),.A2(FE_OFN310_g4336A),.A1(g2257A));
AND2_X1 U_g5148A (.ZN(g5148A),.A2(g4671A),.A1(g1107A));
AND2_X1 U_g9124A (.ZN(g9124A),.A2(FE_OFN325_g18A),.A1(g8881A));
AND2_X1 U_g9324A (.ZN(g9324A),.A2(FE_OFN275_g48A),.A1(g8879A));
AND2_X1 U_g4559A (.ZN(g4559A),.A2(FE_OFN137_g3829A),.A1(g2034A));
AND2_X1 U_g10561A (.ZN(g10561A),.A2(FE_OFN370_g4525A),.A1(g10549A));
AND2_X1 U_g5698A (.ZN(g5698A),.A2(FE_OFN315_g5117A),.A1(g1571A));
AND2_X1 U_g11226A (.ZN(g11226A),.A2(g11060A),.A1(g461A));
AND2_X1 U_g10295A (.ZN(g10295A),.A2(g9995A),.A1(FE_OFN79_g8700A));
AND2_X1 U_g5260A (.ZN(g5260A),.A2(FE_OFN288_g4263A),.A1(g1092A));
AND2_X1 U_g10680A (.ZN(g10680A),.A2(FE_OFN102_g3586A),.A1(g10564A));
AND2_X1 U_g6822A (.ZN(g6822A),.A2(FE_OFN178_g5354A),.A1(g231A));
AND2_X1 U_g4905A (.ZN(g4905A),.A2(g4243A),.A1(g1853A));
AND2_X1 U_g11551A (.ZN(g11551A),.A2(FE_OFN119_g3015A),.A1(g11538A));
AND2_X1 U_g3047A (.ZN(g3047A),.A2(g2306A),.A1(g1227A));
AND2_X1 U_g9849A (.ZN(g9849A),.A2(g9764A),.A1(g293A));
AND2_X1 U_g5279A (.ZN(g5279A),.A2(FE_OFN299_g4457A),.A1(g1766A));
AND2_X1 U_g8404A (.ZN(g8404A),.A2(g8146A),.A1(g686A));
AND2_X1 U_g5720A (.ZN(g5720A),.A2(FE_OFN168_g5361A),.A1(g170A));
AND2_X1 U_g5318A (.ZN(g5318A),.A2(g1857A),.A1(FE_OFN223_g4401A));
AND2_X1 U_g11376A (.ZN(g11376A),.A2(g4285A),.A1(g11318A));
AND2_X1 U_g11297A (.ZN(g11297A),.A2(g11243A),.A1(g4565A));
AND2_X1 U_g9898A (.ZN(g9898A),.A2(g9367A),.A1(g9710A));
OR2_X1 U_g6895A (.ZN(g6895A),.A2(g4875A),.A1(g6776A));
OR2_X1 U_g7189A (.ZN(g7189A),.A2(I9717A),.A1(g6632A));
OR2_X1 U_g9510A (.ZN(g9510A),.A2(g9111A),.A1(FE_OFN44_g9125A));
OR2_X1 U_g7297A (.ZN(g7297A),.A2(g6323A),.A1(g7132A));
OR2_X1 U_g9088A (.ZN(g9088A),.A2(g8233A),.A1(g8927A));
OR2_X1 U_g9923A (.ZN(g9923A),.A2(g9707A),.A1(g9865A));
OR2_X1 U_g6485A (.ZN(g6485A),.A2(g5067A),.A1(g5848A));
OR2_X1 U_g8771A (.ZN(g8771A),.A2(g8652A),.A1(g5483A));
OR2_X1 U_g5813A (.ZN(g5813A),.A2(g4869A),.A1(g5617A));
OR2_X1 U_g7963A (.ZN(g7963A),.A2(g7182A),.A1(FE_OFN334_g7045A));
OR2_X1 U_g10643A (.ZN(g10643A),.A2(g7736A),.A1(g10624A));
OR3_X1 U_g9886A (.ZN(g9886A),.A3(g9759A),.A2(g9592A),.A1(g9607A));
OR3_X1 U_g9951A (.ZN(g9951A),.A3(g9803A),.A2(g9899A),.A1(g9902A));
OR2_X1 U_g11625A (.ZN(g11625A),.A2(g11597A),.A1(g6535A));
OR2_X1 U_g8945A (.ZN(g8945A),.A2(FE_OFN332_g8748A),.A1(g8801A));
OR2_X1 U_g10489A (.ZN(g10489A),.A2(g10367A),.A1(g4456A));
OR2_X1 U_g10559A (.ZN(g10559A),.A2(g10512A),.A1(g4141A));
OR2_X1 U_g10558A (.ZN(g10558A),.A2(g10510A),.A1(g4126A));
OR2_X1 U_g11338A (.ZN(g11338A),.A2(g11178A),.A1(g11283A));
OR2_X1 U_g8435A (.ZN(g8435A),.A2(g8075A),.A1(g8403A));
OR2_X1 U_g10544A (.ZN(g10544A),.A2(g10495A),.A1(g4271A));
OR2_X1 U_g6911A (.ZN(g6911A),.A2(g5681A),.A1(g6342A));
OR2_X1 U_g10865A (.ZN(g10865A),.A2(g10752A),.A1(g5538A));
OR2_X1 U_g3698A (.ZN(g3698A),.A2(g869A),.A1(g3121A));
OR2_X1 U_g8214A (.ZN(g8214A),.A2(g7682A),.A1(g7472A));
OR2_X1 U_g6124A (.ZN(g6124A),.A2(g5188A),.A1(g5181A));
OR2_X1 U_g6469A (.ZN(g6469A),.A2(g4959A),.A1(g5698A));
OR2_X1 U_g5587A (.ZN(g5587A),.A2(g3904A),.A1(g4714A));
OR2_X1 U_g6177A (.ZN(g6177A),.A2(g4712A),.A1(g5444A));
OR2_X1 U_g9891A (.ZN(g9891A),.A2(g9760A),.A1(FE_OFN33_g9454A));
OR2_X1 U_g9913A (.ZN(g9913A),.A2(g9691A),.A1(g9849A));
OR4_X1 U_I5600A (.ZN(I5600A),.A4(g481A),.A3(g486A),.A2(g491A),.A1(g496A));
OR2_X1 U_g11257A (.ZN(g11257A),.A2(g11019A),.A1(g11234A));
OR2_X1 U_g8236A (.ZN(g8236A),.A2(g7680A),.A1(g7526A));
OR2_X1 U_g7385A (.ZN(g7385A),.A2(g6746A),.A1(g7235A));
OR2_X1 U_g6898A (.ZN(g6898A),.A2(g4881A),.A1(g6790A));
OR2_X1 U_g6900A (.ZN(g6900A),.A2(g6246A),.A1(g6787A));
OR2_X1 U_g4264A (.ZN(g4264A),.A2(g4053A),.A1(g4048A));
OR3_X1 U_g9726A (.ZN(g9726A),.A3(g9426A),.A2(g9420A),.A1(g9411A));
OR2_X1 U_g6088A (.ZN(g6088A),.A2(g4522A),.A1(g5260A));
OR2_X1 U_g6923A (.ZN(g6923A),.A2(g5695A),.A1(g6353A));
OR2_X1 U_g8194A (.ZN(g8194A),.A2(g7940A),.A1(g5168A));
OR3_X1 U_g9676A (.ZN(g9676A),.A3(FE_OFN62_g9274A),.A2(FE_OFN72_g9292A),.A1(g9454A));
OR2_X1 U_g11256A (.ZN(g11256A),.A2(g11018A),.A1(g11186A));
OR2_X1 U_g3860A (.ZN(g3860A),.A2(g2167A),.A1(g3107A));
OR2_X1 U_g11280A (.ZN(g11280A),.A2(g11153A),.A1(g11254A));
OR4_X1 U_g9727A (.ZN(g9727A),.A4(I14866A),.A3(g9391A),.A2(g9663A),.A1(g9650A));
OR2_X1 U_g4997A (.ZN(g4997A),.A2(g4584A),.A1(g4581A));
OR2_X1 U_g11624A (.ZN(g11624A),.A2(g11571A),.A1(g11595A));
OR2_X1 U_g11300A (.ZN(g11300A),.A2(g11091A),.A1(g11213A));
OR2_X1 U_g4238A (.ZN(g4238A),.A2(g4007A),.A1(g3999A));
OR2_X1 U_g8814A (.ZN(g8814A),.A2(g8728A),.A1(g7945A));
OR2_X1 U_g10401A (.ZN(g10401A),.A2(g10291A),.A1(g9317A));
OR2_X1 U_g8773A (.ZN(g8773A),.A2(g8653A),.A1(g5491A));
OR2_X1 U_g11231A (.ZN(g11231A),.A2(g11013A),.A1(g11156A));
OR2_X1 U_g10864A (.ZN(g10864A),.A2(g10751A),.A1(g5532A));
OR2_X1 U_g9624A (.ZN(g9624A),.A2(g9313A),.A1(g9316A));
OR3_X1 U_g9953A (.ZN(g9953A),.A3(g9803A),.A2(g9939A),.A1(g9945A));
OR2_X1 U_g6122A (.ZN(g6122A),.A2(g5180A),.A1(g5172A));
OR2_X1 U_g6465A (.ZN(g6465A),.A2(g5041A),.A1(g5825A));
OR2_X1 U_g6934A (.ZN(g6934A),.A2(g5720A),.A1(g6363A));
OR2_X1 U_g7664A (.ZN(g7664A),.A2(FE_OFN350_g3121A),.A1(g6855A));
OR2_X1 U_g7246A (.ZN(g7246A),.A2(g6003A),.A1(g6465A));
OR2_X1 U_g7203A (.ZN(g7203A),.A2(g6058A),.A1(g6640A));
OR2_X1 U_g6096A (.ZN(g6096A),.A2(g4542A),.A1(g5268A));
OR2_X1 U_g9747A (.ZN(g9747A),.A2(g9509A),.A1(g9173A));
OR2_X1 U_g11314A (.ZN(g11314A),.A2(g11102A),.A1(g11224A));
OR2_X1 U_g10733A (.ZN(g10733A),.A2(g10679A),.A1(g5227A));
OR2_X1 U_g8921A (.ZN(g8921A),.A2(g8748A),.A1(g8827A));
OR4_X1 U_I15054A (.ZN(I15054A),.A4(FE_OFN35_g9785A),.A3(FE_OFN61_g9624A),.A2(FE_OFN32_g9454A),.A1(FE_OFN90_I11360A));
OR2_X1 U_g11269A (.ZN(g11269A),.A2(g11031A),.A1(g11196A));
OR2_X1 U_g5555A (.ZN(g5555A),.A2(g4397A),.A1(g4389A));
OR2_X1 U_g11268A (.ZN(g11268A),.A2(g11030A),.A1(g11194A));
OR2_X1 U_g10485A (.ZN(g10485A),.A2(g10363A),.A1(g9317A));
OR2_X1 U_g10555A (.ZN(g10555A),.A2(g10504A),.A1(g4103A));
OR2_X1 U_g6481A (.ZN(g6481A),.A2(g4972A),.A1(g5722A));
OR2_X1 U_g10712A (.ZN(g10712A),.A2(g9097A),.A1(g10662A));
OR2_X1 U_g11335A (.ZN(g11335A),.A2(g11175A),.A1(g11279A));
OR2_X1 U_g8249A (.ZN(g8249A),.A2(g7710A),.A1(g8018A));
OR2_X1 U_g7638A (.ZN(g7638A),.A2(FE_OFN195_g6488A),.A1(g7265A));
OR2_X1 U_g10567A (.ZN(g10567A),.A2(g7378A),.A1(g10514A));
OR2_X1 U_g11487A (.ZN(g11487A),.A2(g11464A),.A1(g6662A));
OR4_X1 U_I15210A (.ZN(I15210A),.A4(g9882A),.A3(g9852A),.A2(g9964A),.A1(g9839A));
OR4_X1 U_I5805A (.ZN(I5805A),.A4(g2088A),.A3(g2096A),.A2(g2099A),.A1(g2102A));
OR2_X1 U_g8941A (.ZN(g8941A),.A2(FE_OFN332_g8748A),.A1(g8796A));
OR2_X1 U_g11443A (.ZN(g11443A),.A2(g11407A),.A1(g7130A));
OR2_X1 U_g4231A (.ZN(g4231A),.A2(g3998A),.A1(g3991A));
OR2_X1 U_g11278A (.ZN(g11278A),.A2(g11150A),.A1(g11253A));
OR2_X1 U_g11286A (.ZN(g11286A),.A2(g11209A),.A1(g10670A));
OR2_X1 U_g8431A (.ZN(g8431A),.A2(g8071A),.A1(g8387A));
OR2_X1 U_g7133A (.ZN(g7133A),.A2(I6273A),.A1(g6616A));
OR2_X1 U_g11306A (.ZN(g11306A),.A2(g11095A),.A1(g11216A));
OR2_X1 U_g8252A (.ZN(g8252A),.A2(g7679A),.A1(g7988A));
OR2_X1 U_g8812A (.ZN(g8812A),.A2(g8724A),.A1(g7939A));
OR2_X1 U_g7846A (.ZN(g7846A),.A2(g7241A),.A1(g7722A));
OR2_X1 U_g3875A (.ZN(g3875A),.A2(g12A),.A1(g3275A));
OR2_X1 U_g5996A (.ZN(g5996A),.A2(g3383A),.A1(g5473A));
OR2_X1 U_g6592A (.ZN(g6592A),.A2(g5882A),.A1(g5100A));
OR2_X1 U_g8286A (.ZN(g8286A),.A2(g7823A),.A1(g8107A));
OR2_X1 U_g10501A (.ZN(g10501A),.A2(g10445A),.A1(g4161A));
OR2_X1 U_g10728A (.ZN(g10728A),.A2(g10642A),.A1(g4973A));
OR2_X1 U_g8270A (.ZN(g8270A),.A2(g3434A),.A1(g7894A));
OR2_X1 U_g7290A (.ZN(g7290A),.A2(g6316A),.A1(g7046A));
OR2_X1 U_g6068A (.ZN(g6068A),.A2(g4497A),.A1(g5220A));
OR2_X1 U_g6468A (.ZN(g6468A),.A2(g4950A),.A1(g5690A));
OR2_X1 U_g11217A (.ZN(g11217A),.A2(g11005A),.A1(g11144A));
OR2_X1 U_g11478A (.ZN(g11478A),.A2(g11455A),.A1(g6532A));
OR4_X2 U_g9536A (.ZN(g9536A),.A4(g9324A),.A3(g9328A),.A2(g9331A),.A1(g9335A));
OR2_X1 U_g5981A (.ZN(g5981A),.A2(g4383A),.A1(g5074A));
OR2_X1 U_g11486A (.ZN(g11486A),.A2(g11463A),.A1(g6654A));
OR2_X1 U_g8377A (.ZN(g8377A),.A2(g7958A),.A1(g8185A));
OR2_X1 U_g8206A (.ZN(g8206A),.A2(g7683A),.A1(g7459A));
OR2_X1 U_g11580A (.ZN(g11580A),.A2(g11544A),.A1(g11413A));
OR2_X1 U_g8287A (.ZN(g8287A),.A2(g7824A),.A1(g8117A));
OR2_X1 U_g11223A (.ZN(g11223A),.A2(g11008A),.A1(g11147A));
OR2_X1 U_g9522A (.ZN(g9522A),.A2(FE_OFN44_g9125A),.A1(g9173A));
OR2_X1 U_g8199A (.ZN(g8199A),.A2(g7444A),.A1(g7902A));
OR2_X1 U_g5802A (.ZN(g5802A),.A2(g4837A),.A1(g5601A));
OR2_X1 U_g11321A (.ZN(g11321A),.A2(g11105A),.A1(g11230A));
OR2_X1 U_g6524A (.ZN(g6524A),.A2(g4996A),.A1(g5746A));
OR2_X1 U_g10664A (.ZN(g10664A),.A2(g10582A),.A1(g10240A));
OR2_X1 U_g7257A (.ZN(g7257A),.A2(g4725A),.A1(g6701A));
OR2_X1 U_g7301A (.ZN(g7301A),.A2(g6327A),.A1(g7140A));
OR2_X1 U_g10484A (.ZN(g10484A),.A2(g10400A),.A1(g9317A));
OR2_X1 U_g10554A (.ZN(g10554A),.A2(g10503A),.A1(g4097A));
OR2_X1 U_g8259A (.ZN(g8259A),.A2(g7719A),.A1(g8028A));
OR2_X1 U_g11334A (.ZN(g11334A),.A2(g11174A),.A1(g11277A));
OR2_X1 U_g8819A (.ZN(g8819A),.A2(g8734A),.A1(g7957A));
OR2_X1 U_g8923A (.ZN(g8923A),.A2(FE_OFN329_g8763A),.A1(g8846A));
OR2_X2 U_g8488A (.ZN(g8488A),.A2(g8390A),.A1(FE_OFN204_g3664A));
OR2_X1 U_g7441A (.ZN(g7441A),.A2(g5867A),.A1(g7271A));
OR2_X1 U_g6026A (.ZN(g6026A),.A2(g3970A),.A1(g5507A));
OR2_X1 U_g10799A (.ZN(g10799A),.A2(g10769A),.A1(g6225A));
OR2_X1 U_g10798A (.ZN(g10798A),.A2(g10768A),.A1(g6217A));
OR2_X1 U_g10805A (.ZN(g10805A),.A2(g10760A),.A1(g10759A));
OR2_X1 U_g10732A (.ZN(g10732A),.A2(g10661A),.A1(g4358A));
OR2_X1 U_g6061A (.ZN(g6061A),.A2(g4A),.A1(g5204A));
OR2_X1 U_g9512A (.ZN(g9512A),.A2(g9125A),.A1(g9151A));
OR2_X1 U_g10013A (.ZN(g10013A),.A2(I15215A),.A1(I15214A));
OR2_X1 U_g8806A (.ZN(g8806A),.A2(g8718A),.A1(g7931A));
OR2_X1 U_g8943A (.ZN(g8943A),.A2(FE_OFN332_g8748A),.A1(g8837A));
OR2_X1 U_g11293A (.ZN(g11293A),.A2(g10818A),.A1(g11211A));
OR2_X1 U_g11265A (.ZN(g11265A),.A2(g11027A),.A1(g11189A));
OR2_X1 U_g8887A (.ZN(g8887A),.A2(FE_OFN329_g8763A),.A1(g8842A));
OR2_X1 U_g5838A (.ZN(g5838A),.A2(g3974A),.A1(g5612A));
OR2_X1 U_g6514A (.ZN(g6514A),.A2(g4992A),.A1(g5738A));
OR2_X1 U_g8322A (.ZN(g8322A),.A2(g6891A),.A1(g8136A));
OR2_X1 U_g8230A (.ZN(g8230A),.A2(g7686A),.A1(g7515A));
OR2_X1 U_g5809A (.ZN(g5809A),.A2(g4865A),.A1(g5611A));
OR2_X1 U_g8433A (.ZN(g8433A),.A2(g8073A),.A1(g8399A));
OR2_X1 U_g11579A (.ZN(g11579A),.A2(g11551A),.A1(g5123A));
OR2_X1 U_g10771A (.ZN(g10771A),.A2(g10684A),.A1(g5533A));
OR2_X1 U_g11615A (.ZN(g11615A),.A2(g11592A),.A1(g11601A));
OR2_X1 U_g9367A (.ZN(g9367A),.A2(g9331A),.A1(g9335A));
OR3_X1 U_g9872A (.ZN(g9872A),.A3(g9759A),.A2(g9594A),.A1(g9617A));
OR2_X1 U_g6522A (.ZN(g6522A),.A2(g4994A),.A1(g5744A));
OR2_X1 U_g8266A (.ZN(g8266A),.A2(g3412A),.A1(g7885A));
OR2_X1 U_g10414A (.ZN(g10414A),.A2(g9291A),.A1(g10300A));
OR2_X1 U_g11275A (.ZN(g11275A),.A2(g11148A),.A1(g11248A));
OR2_X1 U_g11430A (.ZN(g11430A),.A2(g4006A),.A1(g11387A));
OR2_X1 U_g8248A (.ZN(g8248A),.A2(g7707A),.A1(g8014A));
OR2_X1 U_g8815A (.ZN(g8815A),.A2(g8730A),.A1(g7948A));
OR2_X1 U_g7183A (.ZN(g7183A),.A2(I9717A),.A1(g6623A));
OR2_X1 U_g5983A (.ZN(g5983A),.A2(g4392A),.A1(g5084A));
OR2_X1 U_g8154A (.ZN(g8154A),.A2(g6879A),.A1(g7891A));
OR2_X1 U_g6537A (.ZN(g6537A),.A2(g5005A),.A1(g5781A));
OR2_X1 U_g4309A (.ZN(g4309A),.A2(g4079A),.A1(g4069A));
OR2_X1 U_g10725A (.ZN(g10725A),.A2(g10634A),.A1(g4962A));
OR2_X1 U_g6243A (.ZN(g6243A),.A2(g4144A),.A1(g5537A));
OR4_X1 U_I6351A (.ZN(I6351A),.A4(g2372A),.A3(g2380A),.A2(g2389A),.A1(g2405A));
OR3_X1 U_g9519A (.ZN(g9519A),.A3(FE_OFN44_g9125A),.A2(g9151A),.A1(g9173A));
OR2_X1 U_g9740A (.ZN(g9740A),.A2(g9505A),.A1(g9418A));
OR2_X1 U_g8267A (.ZN(g8267A),.A2(g3422A),.A1(g7889A));
OR3_X1 U_g10744A (.ZN(g10744A),.A3(I16427A),.A2(g10668A),.A1(g10381A));
OR2_X1 U_g6542A (.ZN(g6542A),.A2(g5010A),.A1(g5789A));
OR2_X1 U_g7303A (.ZN(g7303A),.A2(g6329A),.A1(g7145A));
OR2_X1 U_g10652A (.ZN(g10652A),.A2(g7743A),.A1(g10627A));
OR2_X1 U_g5036A (.ZN(g5036A),.A2(g4162A),.A1(g4871A));
OR2_X1 U_g7240A (.ZN(g7240A),.A2(g6095A),.A1(g6687A));
OR2_X1 U_g8221A (.ZN(g8221A),.A2(g7688A),.A1(g7496A));
OR2_X1 U_g6902A (.ZN(g6902A),.A2(g4223A),.A1(g6794A));
OR2_X1 U_g10500A (.ZN(g10500A),.A2(g10442A),.A1(g4157A));
OR2_X1 U_g4052A (.ZN(g4052A),.A2(g2515A),.A1(g2862A));
OR4_X1 U_I14858A (.ZN(I14858A),.A4(g9602A),.A3(g9610A),.A2(g9595A),.A1(g9585A));
OR2_X1 U_g6529A (.ZN(g6529A),.A2(g5000A),.A1(g5757A));
OR2_X1 U_g11264A (.ZN(g11264A),.A2(g11026A),.A1(g11188A));
OR4_X1 U_I15209A (.ZN(I15209A),.A4(g9830A),.A3(g9934A),.A2(g9905A),.A1(g8169A));
OR2_X1 U_g8241A (.ZN(g8241A),.A2(g7684A),.A1(g7536A));
OR2_X1 U_g10795A (.ZN(g10795A),.A2(g10764A),.A1(g6199A));
OR2_X1 U_g11607A (.ZN(g11607A),.A2(g11557A),.A1(g11586A));
OR2_X1 U_g8644A (.ZN(g8644A),.A2(g8464A),.A1(g8123A));
OR3_X1 U_g4682A (.ZN(g4682A),.A3(g1570A),.A2(g3348A),.A1(g3563A));
OR2_X1 U_g8818A (.ZN(g8818A),.A2(g8733A),.A1(g7955A));
OR2_X1 U_g2984A (.ZN(g2984A),.A2(g2522A),.A1(g2528A));
OR2_X1 U_g9931A (.ZN(g9931A),.A2(g9900A),.A1(g8931A));
OR2_X1 U_g3414A (.ZN(g3414A),.A2(g2917A),.A1(g2911A));
OR2_X1 U_g9515A (.ZN(g9515A),.A2(g9151A),.A1(g9173A));
OR2_X1 U_g10724A (.ZN(g10724A),.A2(g10672A),.A1(g10312A));
OR2_X1 U_g7294A (.ZN(g7294A),.A2(g6320A),.A1(g7068A));
OR2_X1 U_g5189A (.ZN(g5189A),.A2(FE_OFN292_g3015A),.A1(g4345A));
OR2_X1 U_g8614A (.ZN(g8614A),.A2(g8510A),.A1(g8365A));
OR2_X1 U_g3513A (.ZN(g3513A),.A2(g2180A),.A1(g3118A));
OR2_X1 U_g6909A (.ZN(g6909A),.A2(g5309A),.A1(g6346A));
OR4_X1 U_I5571A (.ZN(I5571A),.A4(g426A),.A3(g386A),.A2(g391A),.A1(g396A));
OR2_X1 U_g4283A (.ZN(g4283A),.A2(g4063A),.A1(g4059A));
OR2_X1 U_g8939A (.ZN(g8939A),.A2(FE_OFN332_g8748A),.A1(g8791A));
OR2_X1 U_g2514A (.ZN(g2514A),.A2(I5600A),.A1(I5599A));
OR2_X1 U_g11327A (.ZN(g11327A),.A2(g11167A),.A1(g11297A));
OR2_X1 U_g8187A (.ZN(g8187A),.A2(g7677A),.A1(g7542A));
OR2_X1 U_g11606A (.ZN(g11606A),.A2(g11556A),.A1(g11585A));
OR2_X1 U_g11303A (.ZN(g11303A),.A2(g11092A),.A1(g11214A));
OR2_X1 U_g5309A (.ZN(g5309A),.A2(g4401A),.A1(FE_OFN204_g3664A));
OR2_X1 U_g8200A (.ZN(g8200A),.A2(g7685A),.A1(g7535A));
OR3_X1 U_g2522A (.ZN(g2522A),.A3(I5629A),.A2(g829A),.A1(g833A));
OR4_X1 U_g2315A (.ZN(g2315A),.A4(I5363A),.A3(g1113A),.A2(g1166A),.A1(g1163A));
OR2_X1 U_g6506A (.ZN(g6506A),.A2(g4989A),.A1(g5731A));
OR2_X1 U_g10649A (.ZN(g10649A),.A2(g7741A),.A1(g10626A));
OR2_X1 U_g8159A (.ZN(g8159A),.A2(g6886A),.A1(g7895A));
OR2_X1 U_g7626A (.ZN(g7626A),.A2(g3440A),.A1(g7060A));
OR2_X1 U_g10770A (.ZN(g10770A),.A2(g10682A),.A1(g5525A));
OR2_X1 U_g11483A (.ZN(g11483A),.A2(g11460A),.A1(g6633A));
OR2_X1 U_g8811A (.ZN(g8811A),.A2(g8722A),.A1(g7935A));
OR3_X1 U_g8642A (.ZN(g8642A),.A3(g8465A),.A2(g31A),.A1(g30A));
OR2_X1 U_g6545A (.ZN(g6545A),.A2(g5025A),.A1(g5795A));
OR2_X1 U_g10767A (.ZN(g10767A),.A2(g10681A),.A1(g5500A));
OR2_X1 U_g11326A (.ZN(g11326A),.A2(g11166A),.A1(g11296A));
OR2_X1 U_g10898A (.ZN(g10898A),.A2(g10777A),.A1(g4220A));
OR2_X1 U_g11252A (.ZN(g11252A),.A2(g10969A),.A1(g11099A));
OR2_X1 U_g10719A (.ZN(g10719A),.A2(g10666A),.A1(g10303A));
OR2_X1 U_g4609A (.ZN(g4609A),.A2(g119A),.A1(g3275A));
OR2_X1 U_g6507A (.ZN(g6507A),.A2(g4990A),.A1(g5732A));
OR2_X1 U_g10718A (.ZN(g10718A),.A2(g10706A),.A1(g6238A));
OR2_X1 U_g10521A (.ZN(g10521A),.A2(I16149A),.A1(I16148A));
OR2_X1 U_g7075A (.ZN(g7075A),.A2(g6530A),.A1(g5104A));
OR2_X1 U_g7292A (.ZN(g7292A),.A2(g6318A),.A1(g7055A));
OR2_X1 U_g10861A (.ZN(g10861A),.A2(g10745A),.A1(g5523A));
OR2_X1 U_g8417A (.ZN(g8417A),.A2(g7721A),.A1(g8246A));
OR2_X1 U_g6515A (.ZN(g6515A),.A2(g4993A),.A1(g5739A));
OR4_X1 U_I14855A (.ZN(I14855A),.A4(g9596A),.A3(g9601A),.A2(g9593A),.A1(g9583A));
OR4_X1 U_I15205A (.ZN(I15205A),.A4(g9878A),.A3(g9850A),.A2(g9963A),.A1(g9838A));
OR4_X1 U_I15051A (.ZN(I15051A),.A4(FE_OFN35_g9785A),.A3(FE_OFN60_g9624A),.A2(g9673A),.A1(FE_OFN90_I11360A));
OR3_X1 U_g9724A (.ZN(g9724A),.A3(g9426A),.A2(g9419A),.A1(g9409A));
OR2_X1 U_g6528A (.ZN(g6528A),.A2(g4999A),.A1(g5756A));
OR2_X1 U_g8823A (.ZN(g8823A),.A2(g8693A),.A1(g8778A));
OR2_X1 U_g7503A (.ZN(g7503A),.A2(g6430A),.A1(g6887A));
OR2_X1 U_g8148A (.ZN(g8148A),.A2(g6872A),.A1(g7884A));
OR2_X1 U_g8649A (.ZN(g8649A),.A2(g3440A),.A1(g8499A));
OR2_X1 U_g3584A (.ZN(g3584A),.A2(g2516A),.A1(g2863A));
OR2_X1 U_g10776A (.ZN(g10776A),.A2(g10758A),.A1(g5544A));
OR3_X1 U_g9680A (.ZN(g9680A),.A3(FE_OFN62_g9274A),.A2(FE_OFN72_g9292A),.A1(FE_OFN32_g9454A));
OR2_X1 U_g10859A (.ZN(g10859A),.A2(g10742A),.A1(g5512A));
OR3_X1 U_I14866A (.ZN(I14866A),.A3(g9619A),.A2(g9609A),.A1(g9590A));
OR2_X1 U_g7299A (.ZN(g7299A),.A2(g6325A),.A1(g7138A));
OR2_X1 U_g10858A (.ZN(g10858A),.A2(g10741A),.A1(g5501A));
OR2_X1 U_g8193A (.ZN(g8193A),.A2(g7937A),.A1(g5145A));
OR3_X1 U_g9511A (.ZN(g9511A),.A3(g9111A),.A2(g9125A),.A1(g9151A));
OR2_X1 U_g7738A (.ZN(g7738A),.A2(g6738A),.A1(g7200A));
OR2_X1 U_g7244A (.ZN(g7244A),.A2(g4720A),.A1(g6699A));
OR2_X1 U_g3425A (.ZN(g3425A),.A2(g2910A),.A1(g2895A));
OR2_X1 U_g7478A (.ZN(g7478A),.A2(g6423A),.A1(g6884A));
OR3_X1 U_g9714A (.ZN(g9714A),.A3(g9654A),.A2(g9366A),.A1(g9664A));
OR2_X1 U_g10025A (.ZN(g10025A),.A2(I15225A),.A1(I15224A));
OR2_X1 U_g6908A (.ZN(g6908A),.A2(g4229A),.A1(g6345A));
OR2_X1 U_g5028A (.ZN(g5028A),.A2(g4128A),.A1(g4836A));
OR2_X1 U_g8253A (.ZN(g8253A),.A2(g7718A),.A1(g8023A));
OR2_X1 U_g8938A (.ZN(g8938A),.A2(FE_OFN332_g8748A),.A1(g8789A));
OR2_X1 U_g8813A (.ZN(g8813A),.A2(g8726A),.A1(g7943A));
OR2_X1 U_g9736A (.ZN(g9736A),.A2(g9423A),.A1(g9430A));
OR2_X1 U_g9968A (.ZN(g9968A),.A2(I15172A),.A1(I15171A));
OR2_X1 U_g8552A (.ZN(g8552A),.A2(g8388A),.A1(g8217A));
OR2_X1 U_g5910A (.ZN(g5910A),.A2(g4341A),.A1(g5023A));
OR2_X1 U_g11249A (.ZN(g11249A),.A2(g11143A),.A1(g6162A));
OR2_X1 U_g11482A (.ZN(g11482A),.A2(g11459A),.A1(g6628A));
OR4_X1 U_g9722A (.ZN(g9722A),.A4(I14855A),.A3(g9391A),.A2(g9643A),.A1(g9612A));
OR4_X1 U_I15204A (.ZN(I15204A),.A4(g9829A),.A3(g9933A),.A2(g9904A),.A1(g8168A));
OR2_X1 U_g7236A (.ZN(g7236A),.A2(g6092A),.A1(g6684A));
OR2_X1 U_g8645A (.ZN(g8645A),.A2(g8469A),.A1(g8127A));
OR2_X1 U_g11647A (.ZN(g11647A),.A2(g11637A),.A1(g6622A));
OR2_X1 U_g6777A (.ZN(g6777A),.A2(g48A),.A1(I9221A));
OR3_X1 U_g9737A (.ZN(g9737A),.A3(g9387A),.A2(g9658A),.A1(g9657A));
OR4_X1 U_I16149A (.ZN(I16149A),.A4(g10467A),.A3(g10468A),.A2(g10470A),.A1(g10472A));
OR2_X1 U_g11233A (.ZN(g11233A),.A2(g10946A),.A1(g11085A));
OR2_X1 U_g8607A (.ZN(g8607A),.A2(g8554A),.A1(g8406A));
OR4_X1 U_I16148A (.ZN(I16148A),.A4(g10474A),.A3(g10476A),.A2(g10384A),.A1(g10386A));
OR2_X1 U_g8158A (.ZN(g8158A),.A2(g6883A),.A1(g7893A));
OR2_X1 U_g5846A (.ZN(g5846A),.A2(g4236A),.A1(g4932A));
OR2_X1 U_g5396A (.ZN(g5396A),.A2(g3684A),.A1(g4481A));
OR2_X1 U_g5803A (.ZN(g5803A),.A2(g3383A),.A1(g5575A));
OR2_X1 U_g11331A (.ZN(g11331A),.A2(g11171A),.A1(g11272A));
OR2_X1 U_g7295A (.ZN(g7295A),.A2(g6321A),.A1(g7071A));
OR2_X1 U_g6541A (.ZN(g6541A),.A2(g5009A),.A1(g5788A));
OR2_X1 U_g8615A (.ZN(g8615A),.A2(g8557A),.A1(g8413A));
OR2_X1 U_g9926A (.ZN(g9926A),.A2(g9715A),.A1(g9868A));
OR2_X1 U_g9754A (.ZN(g9754A),.A2(g9511A),.A1(g9173A));
OR2_X1 U_g8284A (.ZN(g8284A),.A2(g7821A),.A1(g8102A));
OR2_X1 U_g2204A (.ZN(g2204A),.A2(g1394A),.A1(g1393A));
OR2_X1 U_g7471A (.ZN(g7471A),.A2(g6416A),.A1(g6880A));
OR2_X1 U_g7242A (.ZN(g7242A),.A2(g6098A),.A1(g6693A));
OR2_X1 U_g5847A (.ZN(g5847A),.A2(g3987A),.A1(g5626A));
OR2_X1 U_g6901A (.ZN(g6901A),.A2(g6247A),.A1(g6788A));
OR2_X1 U_g8559A (.ZN(g8559A),.A2(g3664A),.A1(g8380A));
OR3_X1 U_g9729A (.ZN(g9729A),.A3(g9387A),.A2(g9357A),.A1(g9618A));
OR2_X1 U_g10860A (.ZN(g10860A),.A2(g10743A),.A1(g5513A));
OR2_X1 U_g9927A (.ZN(g9927A),.A2(g9716A),.A1(g9869A));
OR2_X1 U_g10497A (.ZN(g10497A),.A2(g10396A),.A1(FE_OFN277_g48A));
OR4_X1 U_g9885A (.ZN(g9885A),.A4(g9759A),.A3(g9662A),.A2(g9598A),.A1(g9454A));
OR4_X1 U_g2528A (.ZN(g2528A),.A4(g849A),.A3(g853A),.A2(g857A),.A1(g861A));
OR2_X1 U_g11229A (.ZN(g11229A),.A2(g11012A),.A1(g11154A));
OR2_X1 U_g8973A (.ZN(g8973A),.A2(FE_OFN329_g8763A),.A1(g8821A));
OR2_X1 U_g10658A (.ZN(g10658A),.A2(g7674A),.A1(g10595A));
OR2_X1 U_g10339A (.ZN(g10339A),.A2(g9291A),.A1(g10232A));
OR4_X1 U_I5363A (.ZN(I5363A),.A4(g1160A),.A3(g1157A),.A2(g1153A),.A1(g1149A));
OR2_X1 U_g11310A (.ZN(g11310A),.A2(g11100A),.A1(g11220A));
OR2_X1 U_g6500A (.ZN(g6500A),.A2(g4986A),.A1(g5725A));
OR2_X1 U_g10855A (.ZN(g10855A),.A2(g10736A),.A1(g6075A));
OR2_X1 U_g9916A (.ZN(g9916A),.A2(g9694A),.A1(g9855A));
OR2_X1 U_g10411A (.ZN(g10411A),.A2(g9291A),.A1(g10299A));
OR2_X1 U_g11603A (.ZN(g11603A),.A2(g11553A),.A1(g11582A));
OR4_X1 U_I5357A (.ZN(I5357A),.A4(g1250A),.A3(g1255A),.A2(g1260A),.A1(g1265A));
OR2_X1 U_g6672A (.ZN(g6672A),.A2(g5259A),.A1(g5509A));
OR3_X1 U_g9873A (.ZN(g9873A),.A3(g9758A),.A2(g9599A),.A1(g9623A));
OR2_X1 U_g6523A (.ZN(g6523A),.A2(g4995A),.A1(g5745A));
OR2_X1 U_g10707A (.ZN(g10707A),.A2(g10686A),.A1(g5545A));
OR4_X1 U_I5626A (.ZN(I5626A),.A4(g534A),.A3(g530A),.A2(g525A),.A1(g521A));
OR2_X1 U_g9579A (.ZN(g9579A),.A2(g9030A),.A1(FE_OFN54_g9052A));
OR2_X1 U_g7298A (.ZN(g7298A),.A2(g6324A),.A1(g7136A));
OR2_X1 U_g6551A (.ZN(g6551A),.A2(g5031A),.A1(g5804A));
OR2_X1 U_g6099A (.ZN(g6099A),.A2(g4550A),.A1(g5273A));
OR2_X1 U_g8282A (.ZN(g8282A),.A2(g7819A),.A1(g8101A));
OR2_X1 U_g9917A (.ZN(g9917A),.A2(g9695A),.A1(g9856A));
OR4_X1 U_I15057A (.ZN(I15057A),.A4(FE_OFN35_g9785A),.A3(FE_OFN60_g9624A),.A2(g9680A),.A1(FE_OFN90_I11360A));
OR2_X1 U_g7219A (.ZN(g7219A),.A2(I9717A),.A1(g6661A));
OR2_X1 U_g10019A (.ZN(g10019A),.A2(I15220A),.A1(I15219A));
OR2_X1 U_g5857A (.ZN(g5857A),.A2(g4670A),.A1(g5418A));
OR4_X1 U_g9725A (.ZN(g9725A),.A4(I14862A),.A3(g9391A),.A2(g9659A),.A1(g9642A));
OR2_X1 U_g11298A (.ZN(g11298A),.A2(g11087A),.A1(g11212A));
OR2_X1 U_g10402A (.ZN(g10402A),.A2(g9291A),.A1(g10295A));
OR4_X1 U_g2521A (.ZN(g2521A),.A4(I5626A),.A3(g476A),.A2(g542A),.A1(g538A));
OR2_X1 U_g10866A (.ZN(g10866A),.A2(g10753A),.A1(g5539A));
OR2_X1 U_g6534A (.ZN(g6534A),.A2(g5003A),.A1(g5772A));
OR2_X1 U_g11232A (.ZN(g11232A),.A2(g11015A),.A1(g11158A));
OR3_X1 U_g9706A (.ZN(g9706A),.A3(g9591A),.A2(g9386A),.A1(g9644A));
OR2_X1 U_g10001A (.ZN(g10001A),.A2(I15205A),.A1(I15204A));
OR2_X1 U_g8776A (.ZN(g8776A),.A2(g8655A),.A1(g5510A));
OR2_X1 U_g7225A (.ZN(g7225A),.A2(g6079A),.A1(g6666A));
OR3_X1 U_g9888A (.ZN(g9888A),.A3(g9757A),.A2(g9608A),.A1(g9648A));
OR2_X1 U_g11261A (.ZN(g11261A),.A2(g11023A),.A1(g11238A));
OR3_X1 U_g9956A (.ZN(g9956A),.A3(g9815A),.A2(g9942A),.A1(g9948A));
OR2_X1 U_g10923A (.ZN(g10923A),.A2(g10715A),.A1(g10778A));
OR2_X1 U_g8264A (.ZN(g8264A),.A2(g3912A),.A1(g7879A));
OR2_X1 U_g6513A (.ZN(g6513A),.A2(g4991A),.A1(g5737A));
OR3_X1 U_I14835A (.ZN(I14835A),.A3(g9588A),.A2(g9645A),.A1(g9621A));
OR2_X1 U_g8641A (.ZN(g8641A),.A2(g8463A),.A1(g8120A));
OR3_X1 U_g5361A (.ZN(g5361A),.A3(g126A),.A2(g3348A),.A1(g4316A));
OR2_X1 U_g11316A (.ZN(g11316A),.A2(g11103A),.A1(g11226A));
OR4_X1 U_I16161A (.ZN(I16161A),.A4(g10475A),.A3(g10477A),.A2(g10478A),.A1(g10479A));
OR2_X1 U_g6916A (.ZN(g6916A),.A2(g5687A),.A1(g6348A));
OR2_X1 U_g8777A (.ZN(g8777A),.A2(g8659A),.A1(g5522A));
OR4_X1 U_g2353A (.ZN(g2353A),.A4(g1415A),.A3(g1411A),.A2(g1407A),.A1(g1403A));
OR2_X1 U_g7510A (.ZN(g7510A),.A2(g6730A),.A1(g7186A));
OR3_X1 U_g9957A (.ZN(g9957A),.A3(g9803A),.A2(g9943A),.A1(g9949A));
OR2_X1 U_g2744A (.ZN(g2744A),.A2(I5805A),.A1(I5804A));
OR2_X1 U_g7245A (.ZN(g7245A),.A2(g6102A),.A1(g6696A));
OR2_X1 U_g7291A (.ZN(g7291A),.A2(g6317A),.A1(g7050A));
OR2_X1 U_g8611A (.ZN(g8611A),.A2(g8556A),.A1(g8410A));
OR4_X1 U_I15199A (.ZN(I15199A),.A4(g9828A),.A3(g9932A),.A2(g9903A),.A1(g8167A));
OR2_X1 U_g10550A (.ZN(g10550A),.A2(g10450A),.A1(g4437A));
OR2_X1 U_g11330A (.ZN(g11330A),.A2(g11170A),.A1(g11304A));
OR2_X1 U_g10721A (.ZN(g10721A),.A2(g10669A),.A1(g10306A));
OR2_X1 U_g8153A (.ZN(g8153A),.A2(g6875A),.A1(g7888A));
OR2_X1 U_g10773A (.ZN(g10773A),.A2(g10685A),.A1(g5540A));
OR2_X1 U_g3688A (.ZN(g3688A),.A2(g868A),.A1(g3744A));
OR4_X1 U_I15225A (.ZN(I15225A),.A4(g9881A),.A3(g9859A),.A2(g9967A),.A1(g9842A));
OR2_X1 U_g6042A (.ZN(g6042A),.A2(g3987A),.A1(g5535A));
OR2_X1 U_g10655A (.ZN(g10655A),.A2(g7389A),.A1(g10561A));
OR2_X1 U_g11259A (.ZN(g11259A),.A2(g11021A),.A1(g11236A));
OR2_X1 U_g11225A (.ZN(g11225A),.A2(g11009A),.A1(g11149A));
OR2_X1 U_g5914A (.ZN(g5914A),.A2(g4343A),.A1(g5029A));
OR2_X1 U_g11258A (.ZN(g11258A),.A2(g11020A),.A1(g11235A));
OR2_X1 U_g6054A (.ZN(g6054A),.A2(g4483A),.A1(g5199A));
OR3_X1 U_g9728A (.ZN(g9728A),.A3(g9426A),.A2(g9422A),.A1(g9412A));
OR3_X1 U_g9730A (.ZN(g9730A),.A3(g9423A),.A2(g9425A),.A1(g9414A));
OR2_X1 U_g5820A (.ZN(g5820A),.A2(g3942A),.A1(g5595A));
OR3_X1 U_g8574A (.ZN(g8574A),.A3(g8465A),.A2(I11360A),.A1(g30A));
OR2_X1 U_g11602A (.ZN(g11602A),.A2(g11552A),.A1(g11581A));
OR2_X1 U_g10502A (.ZN(g10502A),.A2(g10503A),.A1(g4169A));
OR2_X1 U_g10557A (.ZN(g10557A),.A2(g10508A),.A1(g4123A));
OR4_X1 U_I15171A (.ZN(I15171A),.A4(g9835A),.A3(g9896A),.A2(g9909A),.A1(g8175A));
OR2_X1 U_g11337A (.ZN(g11337A),.A2(g11177A),.A1(g11282A));
OR2_X1 U_g7465A (.ZN(g7465A),.A2(g6410A),.A1(g6876A));
OR2_X1 U_g8262A (.ZN(g8262A),.A2(g7625A),.A1(g7970A));
OR2_X1 U_g8889A (.ZN(g8889A),.A2(FE_OFN329_g8763A),.A1(g8844A));
OR2_X1 U_g7096A (.ZN(g7096A),.A2(g5911A),.A1(g6544A));
OR2_X1 U_g5995A (.ZN(g5995A),.A2(g5099A),.A1(g5097A));
OR2_X1 U_g8285A (.ZN(g8285A),.A2(g7822A),.A1(g8104A));
OR2_X1 U_g10791A (.ZN(g10791A),.A2(g10762A),.A1(g6186A));
OR2_X1 U_g2499A (.ZN(g2499A),.A2(I5571A),.A1(I5570A));
OR2_X1 U_g6049A (.ZN(g6049A),.A2(g4670A),.A1(g5254A));
OR2_X1 U_g9920A (.ZN(g9920A),.A2(g9701A),.A1(g9860A));
OR2_X1 U_g10556A (.ZN(g10556A),.A2(g10506A),.A1(g4115A));
OR2_X1 U_g8643A (.ZN(g8643A),.A2(g8508A),.A1(g8364A));
OR2_X1 U_g5810A (.ZN(g5810A),.A2(g3912A),.A1(g5588A));
OR2_X1 U_g11336A (.ZN(g11336A),.A2(g11176A),.A1(g11281A));
OR2_X1 U_g8742A (.ZN(g8742A),.A2(g8598A),.A1(g8135A));
OR2_X1 U_g8926A (.ZN(g8926A),.A2(g8763A),.A1(g8848A));
OR2_X1 U_g7218A (.ZN(g7218A),.A2(g6070A),.A1(g6655A));
OR4_X1 U_I15224A (.ZN(I15224A),.A4(g9834A),.A3(g9937A),.A2(g9908A),.A1(g8174A));
OR2_X1 U_g7293A (.ZN(g7293A),.A2(g6319A),.A1(g7063A));
OR2_X1 U_g11288A (.ZN(g11288A),.A2(g11070A),.A1(g11204A));
OR2_X1 U_g10800A (.ZN(g10800A),.A2(g10772A),.A1(g6245A));
OR2_X1 U_g11308A (.ZN(g11308A),.A2(g11098A),.A1(g11218A));
OR2_X1 U_g8269A (.ZN(g8269A),.A2(g3429A),.A1(g7892A));
OR2_X1 U_g10417A (.ZN(g10417A),.A2(g9097A),.A1(g10301A));
OR2_X1 U_g10936A (.ZN(g10936A),.A2(g10808A),.A1(g5170A));
OR2_X1 U_g9388A (.ZN(g9388A),.A2(g9223A),.A1(g9240A));
OR2_X1 U_g6185A (.ZN(g6185A),.A2(g4715A),.A1(g5470A));
OR2_X1 U_g6470A (.ZN(g6470A),.A2(g4960A),.A1(g5699A));
OR2_X1 U_g6897A (.ZN(g6897A),.A2(g6240A),.A1(g6771A));
OR2_X1 U_g8885A (.ZN(g8885A),.A2(FE_OFN329_g8763A),.A1(g8841A));
OR2_X1 U_g11260A (.ZN(g11260A),.A2(g11022A),.A1(g11237A));
OR2_X1 U_g11488A (.ZN(g11488A),.A2(g11465A),.A1(g6671A));
OR2_X1 U_g6105A (.ZN(g6105A),.A2(g4559A),.A1(g5279A));
OR2_X1 U_g10807A (.ZN(g10807A),.A2(g10761A),.A1(g10701A));
OR2_X1 U_g10639A (.ZN(g10639A),.A2(g7734A),.A1(g10623A));
OR2_X1 U_g4556A (.ZN(g4556A),.A2(g1212A),.A1(g3536A));
OR2_X1 U_g8288A (.ZN(g8288A),.A2(g7825A),.A1(g8119A));
OR2_X1 U_g6755A (.ZN(g6755A),.A2(g5479A),.A1(g4934A));
OR3_X1 U_I14862A (.ZN(I14862A),.A3(g9611A),.A2(g9600A),.A1(g9587A));
OR4_X1 U_I16160A (.ZN(I16160A),.A4(g10481A),.A3(g10482A),.A2(g10392A),.A1(g10394A));
OR2_X1 U_g11610A (.ZN(g11610A),.A2(g11560A),.A1(g11589A));
OR4_X1 U_g9711A (.ZN(g9711A),.A4(g9589A),.A3(g9359A),.A2(g9390A),.A1(g9660A));
OR2_X1 U_g6045A (.ZN(g6045A),.A2(g3989A),.A1(g5541A));
OR2_X1 U_g11270A (.ZN(g11270A),.A2(g11032A),.A1(g11198A));
OR2_X1 U_g7258A (.ZN(g7258A),.A2(g5913A),.A1(g6549A));
OR2_X1 U_g6059A (.ZN(g6059A),.A2(g4489A),.A1(g5211A));
OR2_X1 U_g10007A (.ZN(g10007A),.A2(I15210A),.A1(I15209A));
OR2_X1 U_g11267A (.ZN(g11267A),.A2(g11029A),.A1(g11192A));
OR2_X1 U_g11294A (.ZN(g11294A),.A2(g11210A),.A1(g6576A));
OR3_X1 U_g9509A (.ZN(g9509A),.A3(g9111A),.A2(FE_OFN44_g9125A),.A1(g9151A));
OR2_X1 U_g7211A (.ZN(g7211A),.A2(g6067A),.A1(g6647A));
OR2_X1 U_g5404A (.ZN(g5404A),.A2(g3696A),.A1(g4487A));
OR2_X1 U_g4089A (.ZN(g4089A),.A2(I5254A),.A1(g1959A));
OR4_X1 U_I15219A (.ZN(I15219A),.A4(g9833A),.A3(g9936A),.A2(g9907A),.A1(g8172A));
OR2_X1 U_g11219A (.ZN(g11219A),.A2(g11006A),.A1(g11145A));
OR2_X1 U_g6015A (.ZN(g6015A),.A2(g3942A),.A1(g5497A));
OR2_X1 U_g10720A (.ZN(g10720A),.A2(g10667A),.A1(g10304A));
OR2_X1 U_g8265A (.ZN(g8265A),.A2(g4827A),.A1(g7881A));
OR2_X1 U_g5224A (.ZN(g5224A),.A2(g3512A),.A1(g4360A));
OR3_X1 U_g9700A (.ZN(g9700A),.A3(I14827A),.A2(g9667A),.A1(g9358A));
OR2_X1 U_g7106A (.ZN(g7106A),.A2(g5917A),.A1(g6554A));
OR2_X1 U_g8770A (.ZN(g8770A),.A2(g8651A),.A1(g5476A));
OR2_X1 U_g11201A (.ZN(g11201A),.A2(g11011A),.A1(g11152A));
OR3_X1 U_g9950A (.ZN(g9950A),.A3(g9803A),.A2(g9898A),.A1(g9901A));
OR4_X1 U_g9723A (.ZN(g9723A),.A4(I14858A),.A3(g9391A),.A2(g9652A),.A1(g9620A));
OR2_X1 U_g2309A (.ZN(g2309A),.A2(I5358A),.A1(I5357A));
OR2_X1 U_g11266A (.ZN(g11266A),.A2(g11028A),.A1(g11190A));
OR2_X1 U_g10727A (.ZN(g10727A),.A2(g10638A),.A1(g4969A));
OR2_X1 U_g10863A (.ZN(g10863A),.A2(g10750A),.A1(g5531A));
OR2_X1 U_g8429A (.ZN(g8429A),.A2(g8069A),.A1(g8385A));
OR2_X1 U_g9751A (.ZN(g9751A),.A2(g9510A),.A1(g9515A));
OR2_X1 U_g8281A (.ZN(g8281A),.A2(g7818A),.A1(g8097A));
OR2_X1 U_g6910A (.ZN(g6910A),.A2(g5680A),.A1(g6341A));
OR2_X1 U_g8639A (.ZN(g8639A),.A2(g8462A),.A1(g8118A));
OR3_X1 U_g9673A (.ZN(g9673A),.A3(g9274A),.A2(FE_OFN72_g9292A),.A1(g9454A));
OR2_X1 U_g11285A (.ZN(g11285A),.A2(g11161A),.A1(g11255A));
OR2_X1 U_g11305A (.ZN(g11305A),.A2(g11093A),.A1(g11215A));
OR4_X1 U_I15177A (.ZN(I15177A),.A4(g9876A),.A3(g9863A),.A2(g9960A),.A1(g9844A));
OR3_X1 U_g9734A (.ZN(g9734A),.A3(g9426A),.A2(g9428A),.A1(g9415A));
OR3_X1 U_I14827A (.ZN(I14827A),.A3(g9584A),.A2(g9614A),.A1(g9603A));
OR2_X1 U_g5824A (.ZN(g5824A),.A2(g4839A),.A1(g5602A));
OR2_X1 U_g8715A (.ZN(g8715A),.A2(g8687A),.A1(g8416A));
OR2_X1 U_g5762A (.ZN(g5762A),.A2(g5186A),.A1(g5178A));
OR2_X1 U_g6538A (.ZN(g6538A),.A2(g5006A),.A1(g5782A));
OR2_X1 U_g5590A (.ZN(g5590A),.A2(g4723A),.A1(g4718A));
OR2_X1 U_g10726A (.ZN(g10726A),.A2(g10673A),.A1(g10316A));
OR2_X1 U_g3120A (.ZN(g3120A),.A2(I6351A),.A1(I6350A));
OR3_X2 U_g4640A (.ZN(g4640A),.A3(g1527A),.A2(g3563A),.A1(g3348A));
OR2_X1 U_g6093A (.ZN(g6093A),.A2(g4534A),.A1(g5264A));
OR2_X1 U_g8162A (.ZN(g8162A),.A2(g6889A),.A1(g7898A));
OR2_X1 U_g8268A (.ZN(g8268A),.A2(g7613A),.A1(g7962A));
OR2_X1 U_g9569A (.ZN(g9569A),.A2(FE_OFN49_g9030A),.A1(FE_OFN54_g9052A));
OR2_X1 U_g11485A (.ZN(g11485A),.A2(g11462A),.A1(g6646A));
OR2_X1 U_g10797A (.ZN(g10797A),.A2(g10766A),.A1(g6206A));
OR3_X1 U_I14779A (.ZN(I14779A),.A3(g9192A),.A2(g9205A),.A1(g8995A));
OR2_X1 U_g10408A (.ZN(g10408A),.A2(g9097A),.A1(g10298A));
OR2_X1 U_g10635A (.ZN(g10635A),.A2(g7732A),.A1(g10622A));
OR2_X1 U_g2305A (.ZN(g2305A),.A2(I5352A),.A1(I5351A));
OR4_X1 U_I15176A (.ZN(I15176A),.A4(g9836A),.A3(g9897A),.A2(g9908A),.A1(g8176A));
OR2_X1 U_g3435A (.ZN(g3435A),.A2(g2950A),.A1(g2945A));
OR2_X1 U_g9924A (.ZN(g9924A),.A2(g9709A),.A1(g9866A));
OR2_X1 U_g10711A (.ZN(g10711A),.A2(g10690A),.A1(g5547A));
OR2_X1 U_g5814A (.ZN(g5814A),.A2(g4827A),.A1(g5591A));
OR2_X1 U_g5038A (.ZN(g5038A),.A2(g4884A),.A1(g4878A));
OR4_X1 U_I15215A (.ZN(I15215A),.A4(g9879A),.A3(g9854A),.A2(g9965A),.A1(g9840A));
OR2_X1 U_g8226A (.ZN(g8226A),.A2(g7681A),.A1(g7504A));
OR2_X1 U_g7367A (.ZN(g7367A),.A2(g6744A),.A1(g7224A));
OR2_X1 U_g7457A (.ZN(g7457A),.A2(g6404A),.A1(g6873A));
OR2_X1 U_g5229A (.ZN(g5229A),.A2(g3516A),.A1(g4364A));
OR2_X1 U_g5993A (.ZN(g5993A),.A2(g4400A),.A1(g5090A));
OR2_X1 U_g8283A (.ZN(g8283A),.A2(g7820A),.A1(g8098A));
OR2_X1 U_g7971A (.ZN(g7971A),.A2(g7549A),.A1(g5110A));
OR2_X1 U_g8602A (.ZN(g8602A),.A2(g8550A),.A1(g8401A));
OR2_X1 U_g8920A (.ZN(g8920A),.A2(FE_OFN329_g8763A),.A1(g8845A));
OR2_X1 U_g10663A (.ZN(g10663A),.A2(g10581A),.A1(g10237A));
OR2_X1 U_g6074A (.ZN(g6074A),.A2(g1A),.A1(g5349A));
OR2_X1 U_g8261A (.ZN(g8261A),.A2(g3383A),.A1(g7876A));
OR2_X1 U_g10862A (.ZN(g10862A),.A2(g10746A),.A1(g5524A));
OR2_X1 U_g5837A (.ZN(g5837A),.A2(g4224A),.A1(g5640A));
OR2_X1 U_g11333A (.ZN(g11333A),.A2(g11173A),.A1(g11274A));
OR2_X1 U_g6080A (.ZN(g6080A),.A2(g4512A),.A1(g5249A));
OR2_X1 U_g6480A (.ZN(g6480A),.A2(g4971A),.A1(g5721A));
OR2_X1 U_g7740A (.ZN(g7740A),.A2(g6741A),.A1(g7209A));
OR2_X2 U_g10702A (.ZN(g10702A),.A2(g2984A),.A1(g10562A));
OR3_X1 U_g9697A (.ZN(g9697A),.A3(I14822A),.A2(g9606A),.A1(g9665A));
OR2_X1 U_g8203A (.ZN(g8203A),.A2(g7696A),.A1(g7453A));
OR2_X1 U_g9914A (.ZN(g9914A),.A2(g9692A),.A1(g9851A));
OR2_X1 U_g10564A (.ZN(g10564A),.A2(g7368A),.A1(g10560A));
OR2_X1 U_g11484A (.ZN(g11484A),.A2(g11461A),.A1(g6639A));
OR2_X1 U_g5842A (.ZN(g5842A),.A2(g3979A),.A1(g5618A));
OR4_X1 U_I15200A (.ZN(I15200A),.A4(g9880A),.A3(g9848A),.A2(g9962A),.A1(g9837A));
OR2_X1 U_g11609A (.ZN(g11609A),.A2(g11559A),.A1(g11588A));
OR2_X1 U_g8940A (.ZN(g8940A),.A2(FE_OFN332_g8748A),.A1(g8793A));
OR2_X1 U_g11312A (.ZN(g11312A),.A2(g11101A),.A1(g11222A));
OR2_X1 U_g11608A (.ZN(g11608A),.A2(g11558A),.A1(g11587A));
OR2_X1 U_g6000A (.ZN(g6000A),.A2(g3912A),.A1(g5480A));
OR2_X1 U_g8428A (.ZN(g8428A),.A2(g8068A),.A1(g8382A));
OR2_X1 U_g8430A (.ZN(g8430A),.A2(g8070A),.A1(g8386A));
OR2_X1 U_g9922A (.ZN(g9922A),.A2(g9705A),.A1(g9864A));
OR2_X1 U_g8247A (.ZN(g8247A),.A2(g7704A),.A1(g8010A));
OR2_X1 U_g3438A (.ZN(g3438A),.A2(g2944A),.A1(g2939A));
OR4_X1 U_I5576A (.ZN(I5576A),.A4(g444A),.A3(g440A),.A2(g435A),.A1(g431A));
OR2_X1 U_g6924A (.ZN(g6924A),.A2(g4261A),.A1(g6362A));
OR2_X1 U_g5405A (.ZN(g5405A),.A2(FE_OFN221_g3440A),.A1(g4476A));
OR2_X1 U_g8638A (.ZN(g8638A),.A2(g8461A),.A1(g8108A));
OR2_X1 U_g8609A (.ZN(g8609A),.A2(g8555A),.A1(g8408A));
OR2_X1 U_g9995A (.ZN(g9995A),.A2(I15200A),.A1(I15199A));
OR2_X1 U_g8883A (.ZN(g8883A),.A2(FE_OFN329_g8763A),.A1(g8838A));
OR4_X1 U_I15214A (.ZN(I15214A),.A4(g9831A),.A3(g9935A),.A2(g9906A),.A1(g8170A));
OR3_X1 U_g2538A (.ZN(g2538A),.A3(I5649A),.A2(g1458A),.A1(g1466A));
OR2_X1 U_g11329A (.ZN(g11329A),.A2(g11169A),.A1(g11302A));
OR2_X1 U_g4255A (.ZN(g4255A),.A2(g4047A),.A1(g4009A));
OR2_X1 U_g11328A (.ZN(g11328A),.A2(g11168A),.A1(g11299A));
OR3_X1 U_g9704A (.ZN(g9704A),.A3(I14835A),.A2(g9605A),.A1(g9385A));
OR4_X1 U_I5352A (.ZN(I5352A),.A4(g1117A),.A3(g1121A),.A2(g1125A),.A1(g1129A));
OR2_X1 U_g8774A (.ZN(g8774A),.A2(g8654A),.A1(g5499A));
OR3_X1 U_g9954A (.ZN(g9954A),.A3(g9803A),.A2(g9940A),.A1(g9946A));
OR2_X1 U_g10405A (.ZN(g10405A),.A2(g9291A),.A1(g10297A));
OR2_X1 U_g9363A (.ZN(g9363A),.A2(g9192A),.A1(g9205A));
OR2_X1 U_g5849A (.ZN(g5849A),.A2(g4144A),.A1(g4949A));
OR4_X1 U_I5599A (.ZN(I5599A),.A4(g501A),.A3(g506A),.A2(g511A),.A1(g516A));
OR2_X1 U_g7204A (.ZN(g7204A),.A2(I9717A),.A1(g6645A));
OR2_X1 U_g7300A (.ZN(g7300A),.A2(g6326A),.A1(g7139A));
OR2_X1 U_g4293A (.ZN(g4293A),.A2(g4068A),.A1(g4064A));
OR2_X1 U_g9912A (.ZN(g9912A),.A2(g9690A),.A1(g9847A));
OR2_X1 U_g6533A (.ZN(g6533A),.A2(g5002A),.A1(g5771A));
OR2_X1 U_g8816A (.ZN(g8816A),.A2(g8731A),.A1(g7951A));
OR2_X1 U_g9929A (.ZN(g9929A),.A2(g9718A),.A1(g9871A));
OR2_X1 U_g5819A (.ZN(g5819A),.A2(g4876A),.A1(g5625A));
OR3_X1 U_I14831A (.ZN(I14831A),.A3(g9586A),.A2(g9622A),.A1(g9613A));
OR2_X1 U_g5852A (.ZN(g5852A),.A2(g3989A),.A1(g5632A));
OR2_X1 U_g8263A (.ZN(g8263A),.A2(g7720A),.A1(g8032A));
OR2_X1 U_g3431A (.ZN(g3431A),.A2(g2957A),.A1(g2951A));
OR2_X1 U_g8631A (.ZN(g8631A),.A2(g7449A),.A1(g8474A));
OR2_X1 U_g6922A (.ZN(g6922A),.A2(g5694A),.A1(g6352A));
OR2_X1 U_g8817A (.ZN(g8817A),.A2(g8732A),.A1(g7954A));
OR4_X1 U_g9735A (.ZN(g9735A),.A4(g9387A),.A3(g9384A),.A2(g9651A),.A1(g9649A));
OR2_X1 U_g8605A (.ZN(g8605A),.A2(g8553A),.A1(g8404A));
OR2_X1 U_g11263A (.ZN(g11263A),.A2(g11025A),.A1(g11187A));
OR2_X1 U_g6739A (.ZN(g6739A),.A2(g5780A),.A1(g5769A));
OR2_X1 U_g11332A (.ZN(g11332A),.A2(g11172A),.A1(g11273A));
OR2_X1 U_g7143A (.ZN(g7143A),.A2(I9717A),.A1(g6619A));
OR2_X1 U_g6479A (.ZN(g6479A),.A2(g4968A),.A1(g5707A));
OR4_X1 U_I15048A (.ZN(I15048A),.A4(FE_OFN35_g9785A),.A3(FE_OFN61_g9624A),.A2(g9680A),.A1(FE_OFN90_I11360A));
OR2_X1 U_g6501A (.ZN(g6501A),.A2(g4987A),.A1(g5726A));
OR3_X1 U_g9702A (.ZN(g9702A),.A3(I14831A),.A2(g9647A),.A1(g9365A));
OR2_X1 U_g11221A (.ZN(g11221A),.A2(g11007A),.A1(g11146A));
OR3_X1 U_g9952A (.ZN(g9952A),.A3(g9815A),.A2(g9938A),.A1(g9944A));
OR2_X1 U_g11613A (.ZN(g11613A),.A2(g11591A),.A1(g11600A));
OR2_X1 U_g7621A (.ZN(g7621A),.A2(g6994A),.A1(g5108A));
OR2_X1 U_g3399A (.ZN(g3399A),.A2(g2940A),.A1(g2918A));
OR2_X1 U_g11605A (.ZN(g11605A),.A2(g11555A),.A1(g11584A));
OR2_X1 U_g4274A (.ZN(g4274A),.A2(g4058A),.A1(g4054A));
OR3_X1 U_I14602A (.ZN(I14602A),.A3(g9192A),.A2(FE_OFN42_g9205A),.A1(g8995A));
OR4_X1 U_I15033A (.ZN(I15033A),.A4(FE_OFN35_g9785A),.A3(FE_OFN61_g9624A),.A2(FE_OFN33_g9454A),.A1(FE_OFN90_I11360A));
OR2_X1 U_g10717A (.ZN(g10717A),.A2(g10705A),.A1(g6235A));
OR3_X1 U_I5629A (.ZN(I5629A),.A3(g837A),.A2(g841A),.A1(g845A));
OR2_X1 U_g9925A (.ZN(g9925A),.A2(g9712A),.A1(g9867A));
OR2_X1 U_g3819A (.ZN(g3819A),.A2(g9A),.A1(g3275A));
OR2_X1 U_g6912A (.ZN(g6912A),.A2(g4235A),.A1(g6350A));
OR2_X1 U_g10723A (.ZN(g10723A),.A2(g10633A),.A1(g4952A));
OR2_X1 U_g6929A (.ZN(g6929A),.A2(g5704A),.A1(g6360A));
OR2_X1 U_g10646A (.ZN(g10646A),.A2(g7739A),.A1(g10625A));
OR2_X1 U_g9516A (.ZN(g9516A),.A2(FE_OFN44_g9125A),.A1(FE_OFN47_g9151A));
OR2_X1 U_g6626A (.ZN(g6626A),.A2(g123A),.A1(g5934A));
OR4_X1 U_I6350A (.ZN(I6350A),.A4(g2419A),.A3(g2433A),.A2(g2437A),.A1(g2445A));
OR2_X1 U_g11325A (.ZN(g11325A),.A2(g11165A),.A1(g11295A));
OR4_X1 U_I5366A (.ZN(I5366A),.A4(g1296A),.A3(g1292A),.A2(g1284A),.A1(g1280A));
OR3_X1 U_I5649A (.ZN(I5649A),.A3(g1482A),.A2(g1486A),.A1(g1499A));
OR2_X1 U_g6894A (.ZN(g6894A),.A2(g4868A),.A1(g6763A));
OR3_X1 U_g9738A (.ZN(g9738A),.A3(g9506A),.A2(g9447A),.A1(g9417A));
OR2_X1 U_g8383A (.ZN(g8383A),.A2(g5051A),.A1(g8163A));
OR2_X1 U_g8779A (.ZN(g8779A),.A2(g8663A),.A1(g5530A));
OR2_X1 U_g8161A (.ZN(g8161A),.A2(g7185A),.A1(g8005A));
OR2_X2 U_g8451A (.ZN(g8451A),.A2(g8366A),.A1(FE_OFN221_g3440A));
OR2_X1 U_g9915A (.ZN(g9915A),.A2(g9693A),.A1(g9853A));
OR4_X1 U_g2316A (.ZN(g2316A),.A4(I5366A),.A3(g1270A),.A2(g1304A),.A1(g1300A));
OR2_X1 U_g5576A (.ZN(g5576A),.A2(FE_OFN204_g3664A),.A1(g4675A));
OR2_X1 U_g10857A (.ZN(g10857A),.A2(g10738A),.A1(g6090A));
OR2_X1 U_g10793A (.ZN(g10793A),.A2(g10763A),.A1(g6194A));
OR2_X1 U_g7511A (.ZN(g7511A),.A2(g6438A),.A1(g6890A));
OR2_X1 U_g8944A (.ZN(g8944A),.A2(FE_OFN332_g8748A),.A1(g8799A));
OR2_X1 U_g10765A (.ZN(g10765A),.A2(g10680A),.A1(g5492A));
OR2_X1 U_g10549A (.ZN(g10549A),.A2(g10451A),.A1(g4271A));
OR2_X1 U_g7092A (.ZN(g7092A),.A2(g5902A),.A1(g6540A));
OR2_X1 U_g11604A (.ZN(g11604A),.A2(g11554A),.A1(g11583A));
OR2_X1 U_g8434A (.ZN(g8434A),.A2(g8074A),.A1(g8400A));
OR2_X1 U_g6546A (.ZN(g6546A),.A2(g5026A),.A1(g5796A));
OR2_X1 U_g3354A (.ZN(g3354A),.A2(g1216A),.A1(g3121A));
OR2_X1 U_g9928A (.ZN(g9928A),.A2(g9717A),.A1(g9870A));
OR2_X1 U_g11262A (.ZN(g11262A),.A2(g11024A),.A1(g11240A));
OR4_X1 U_g9785A (.ZN(g9785A),.A4(g9363A),.A3(g9388A),.A2(g8995A),.A1(g9010A));
OR2_X1 U_g5867A (.ZN(g5867A),.A2(g4921A),.A1(FE_OFN221_g3440A));
OR2_X1 U_g8210A (.ZN(g8210A),.A2(g7692A),.A1(g7466A));
OR2_X1 U_g10533A (.ZN(g10533A),.A2(g10449A),.A1(g4437A));
OR2_X1 U_g9563A (.ZN(g9563A),.A2(g9030A),.A1(FE_OFN56_g9052A));
OR2_X1 U_g6906A (.ZN(g6906A),.A2(g5674A),.A1(g6791A));
OR2_X1 U_g7375A (.ZN(g7375A),.A2(g6745A),.A1(g7230A));
OR2_X1 U_g7651A (.ZN(g7651A),.A2(FE_OFN350_g3121A),.A1(g7135A));
OR4_X1 U_I5570A (.ZN(I5570A),.A4(g401A),.A3(g406A),.A2(g411A),.A1(g416A));
OR3_X1 U_g9731A (.ZN(g9731A),.A3(g9387A),.A2(g9364A),.A1(g9641A));
OR2_X1 U_g11247A (.ZN(g11247A),.A2(g10949A),.A1(g11097A));
OR4_X1 U_I15045A (.ZN(I15045A),.A4(FE_OFN35_g9785A),.A3(FE_OFN61_g9624A),.A2(g9676A),.A1(FE_OFN90_I11360A));
OR2_X1 U_g10856A (.ZN(g10856A),.A2(g10737A),.A1(g6083A));
OR2_X1 U_g7184A (.ZN(g7184A),.A2(g6047A),.A1(g6625A));
OR2_X1 U_g11612A (.ZN(g11612A),.A2(g11590A),.A1(g11599A));
OR2_X1 U_g7384A (.ZN(g7384A),.A2(g6618A),.A1(g7088A));
OR2_X1 U_g11324A (.ZN(g11324A),.A2(g11164A),.A1(g11271A));
OR2_X1 U_g8922A (.ZN(g8922A),.A2(FE_OFN329_g8763A),.A1(g8822A));
OR4_X1 U_I5358A (.ZN(I5358A),.A4(g1275A),.A3(g1235A),.A2(g1240A),.A1(g1245A));
OR3_X1 U_g9955A (.ZN(g9955A),.A3(g9803A),.A2(g9941A),.A1(g9947A));
OR4_X1 U_g2501A (.ZN(g2501A),.A4(I5576A),.A3(g421A),.A2(g452A),.A1(g448A));
OR2_X1 U_g7231A (.ZN(g7231A),.A2(g6087A),.A1(g6673A));
OR2_X1 U_g6078A (.ZN(g6078A),.A2(g5256A),.A1(g4503A));
OR2_X1 U_g6478A (.ZN(g6478A),.A2(g4967A),.A1(g5706A));
OR2_X1 U_g6907A (.ZN(g6907A),.A2(g5675A),.A1(g6792A));
OR2_X1 U_g6035A (.ZN(g6035A),.A2(g3974A),.A1(g5518A));
OR2_X1 U_g8937A (.ZN(g8937A),.A2(FE_OFN332_g8748A),.A1(g8786A));
OR2_X1 U_g7742A (.ZN(g7742A),.A2(g6743A),.A1(g7217A));
OR2_X1 U_g10722A (.ZN(g10722A),.A2(g10671A),.A1(g10308A));
OR2_X1 U_g9918A (.ZN(g9918A),.A2(g9698A),.A1(g9858A));
OR2_X1 U_g5403A (.ZN(g5403A),.A2(g3695A),.A1(g4486A));
OR2_X1 U_g7926A (.ZN(g7926A),.A2(g6892A),.A1(g7435A));
OR2_X1 U_g6915A (.ZN(g6915A),.A2(g5686A),.A1(g6347A));
OR2_X1 U_g5841A (.ZN(g5841A),.A2(g4230A),.A1(g4914A));
OR4_X1 U_I15220A (.ZN(I15220A),.A4(g9877A),.A3(g9857A),.A2(g9966A),.A1(g9841A));
OR2_X1 U_g10529A (.ZN(g10529A),.A2(I16161A),.A1(I16160A));
OR2_X1 U_g11246A (.ZN(g11246A),.A2(g10948A),.A1(g11094A));
OR2_X1 U_g6002A (.ZN(g6002A),.A2(g4827A),.A1(g5489A));
OR2_X1 U_g7712A (.ZN(g7712A),.A2(FE_OFN350_g3121A),.A1(g7125A));
OR2_X1 U_g8810A (.ZN(g8810A),.A2(g8720A),.A1(g7933A));
OR2_X1 U_g9921A (.ZN(g9921A),.A2(g9703A),.A1(g9862A));
OR2_X1 U_g8432A (.ZN(g8432A),.A2(g8072A),.A1(g8389A));
OR4_X1 U_I15172A (.ZN(I15172A),.A4(g9874A),.A3(g9861A),.A2(g9959A),.A1(g9843A));
OR3_X1 U_I14822A (.ZN(I14822A),.A3(g9582A),.A2(g9604A),.A1(g9597A));
OR2_X1 U_g6928A (.ZN(g6928A),.A2(g5703A),.A1(g6359A));
OR2_X1 U_g8157A (.ZN(g8157A),.A2(g7623A),.A1(FE_OFN192_g6488A));
OR2_X1 U_g6930A (.ZN(g6930A),.A2(g4269A),.A1(g6364A));
OR2_X1 U_g7660A (.ZN(g7660A),.A2(g5867A),.A1(g7059A));
OR2_X1 U_g6899A (.ZN(g6899A),.A2(g32A),.A1(g6463A));
OR2_X1 U_g9392A (.ZN(g9392A),.A2(g9324A),.A1(g9328A));
OR2_X1 U_g11318A (.ZN(g11318A),.A2(g11104A),.A1(g11228A));
OR3_X1 U_I16427A (.ZN(I16427A),.A3(g10382A),.A2(g10383A),.A1(g10683A));
OR2_X1 U_g11227A (.ZN(g11227A),.A2(g11010A),.A1(g11151A));
OR2_X1 U_g11058A (.ZN(g11058A),.A2(g5280A),.A1(g10933A));
OR4_X1 U_I5351A (.ZN(I5351A),.A4(g1133A),.A3(g1137A),.A2(g1141A),.A1(g1145A));
OR3_X1 U_g9708A (.ZN(g9708A),.A3(g9646A),.A2(g9389A),.A1(g9653A));
OR2_X1 U_g6071A (.ZN(g6071A),.A2(g4505A),.A1(g5228A));
OR2_X1 U_g9911A (.ZN(g9911A),.A2(g9689A),.A1(g9846A));
OR2_X1 U_g7102A (.ZN(g7102A),.A2(g5915A),.A1(g6550A));
OR2_X1 U_g7302A (.ZN(g7302A),.A2(g6328A),.A1(g7141A));
OR2_X1 U_g6038A (.ZN(g6038A),.A2(g3979A),.A1(g5528A));
OR2_X1 U_g4239A (.ZN(g4239A),.A2(g4008A),.A1(g4000A));
OR2_X1 U_g8646A (.ZN(g8646A),.A2(g8547A),.A1(g8224A));
OR2_X1 U_g9974A (.ZN(g9974A),.A2(I15177A),.A1(I15176A));
OR2_X1 U_g5823A (.ZN(g5823A),.A2(g4882A),.A1(g5631A));
OR2_X1 U_g6918A (.ZN(g6918A),.A2(g4252A),.A1(g6358A));
OR2_X1 U_g7265A (.ZN(g7265A),.A2(g6204A),.A1(g6756A));
OR4_X1 U_I5804A (.ZN(I5804A),.A4(g2104A),.A3(g2106A),.A2(g2109A),.A1(g2111A));
OR2_X1 U_g5851A (.ZN(g5851A),.A2(g4253A),.A1(g4941A));
OR2_X1 U_g11481A (.ZN(g11481A),.A2(g11458A),.A1(g6624A));
OR2_X1 U_g10336A (.ZN(g10336A),.A2(g9097A),.A1(g10230A));
OR2_X1 U_g7296A (.ZN(g7296A),.A2(g6322A),.A1(g7131A));
OR2_X1 U_g4300A (.ZN(g4300A),.A2(g1212A),.A1(g3546A));
OR2_X1 U_g8647A (.ZN(g8647A),.A2(g8470A),.A1(g8130A));
NAND2_X1 U_g8546A (.ZN(g8546A),.A2(g8390A),.A1(g3983A));
NAND2_X1 U_g2516A (.ZN(g2516A),.A2(I5613A),.A1(I5612A));
NAND2_X1 U_g2987A (.ZN(g2987A),.A2(g883A),.A1(g2481A));
NAND2_X1 U_I5593A (.ZN(I5593A),.A2(I5591A),.A1(g1703A));
NAND2_X1 U_g8970A (.ZN(g8970A),.A2(g8839A),.A1(g5548A));
NAND2_X1 U_I10519A (.ZN(I10519A),.A2(g822A),.A1(g6231A));
NAND2_X1 U_I11279A (.ZN(I11279A),.A2(I11278A),.A1(g305A));
NAND4_X1 U_g7990A (.ZN(g7990A),.A4(g7550A),.A3(g7562A),.A2(FE_OFN80_g2175A),.A1(FE_OFN88_g2178A));
NAND2_X1 U_I11278A (.ZN(I11278A),.A2(g6485A),.A1(g305A));
NAND2_X1 U_g3978A (.ZN(g3978A),.A2(g1822A),.A1(g3207A));
NAND2_X1 U_I5264A (.ZN(I5264A),.A2(I5263A),.A1(g456A));
NAND2_X1 U_I8640A (.ZN(I8640A),.A2(g516A),.A1(g4278A));
NAND2_X1 U_I6761A (.ZN(I6761A),.A2(I6760A),.A1(g2943A));
NAND2_X1 U_I17400A (.ZN(I17400A),.A2(g11416A),.A1(g11418A));
NAND2_X1 U_I5450A (.ZN(I5450A),.A2(I5449A),.A1(g1235A));
NAND2_X1 U_I16060A (.ZN(I16060A),.A2(I16058A),.A1(g10441A));
NAND2_X1 U_I6746A (.ZN(I6746A),.A2(g1453A),.A1(g2938A));
NAND2_X1 U_I11975A (.ZN(I11975A),.A2(I11973A),.A1(g1462A));
NAND2_X1 U_I12136A (.ZN(I12136A),.A2(g131A),.A1(g6038A));
NAND2_X1 U_I11937A (.ZN(I11937A),.A2(I11935A),.A1(g1458A));
NAND2_X1 U_g2959A (.ZN(g2959A),.A2(I6168A),.A1(I6167A));
NAND2_X1 U_I5878A (.ZN(I5878A),.A2(g2115A),.A1(g2120A));
NAND2_X1 U_g2517A (.ZN(g2517A),.A2(I5620A),.A1(I5619A));
NAND2_X1 U_g5552A (.ZN(g5552A),.A2(FE_OFN223_g4401A),.A1(g4777A));
NAND2_X1 U_I6468A (.ZN(I6468A),.A2(I6467A),.A1(g23A));
NAND2_X1 U_I8796A (.ZN(I8796A),.A2(I8795A),.A1(g4672A));
NAND2_X1 U_g10392A (.ZN(g10392A),.A2(I15892A),.A1(I15891A));
NAND2_X1 U_I5611A (.ZN(I5611A),.A2(g1284A),.A1(g1280A));
NAND2_X1 U_g8738A (.ZN(g8738A),.A2(FE_OFN200_g4921A),.A1(g8688A));
NAND2_X1 U_I6716A (.ZN(I6716A),.A2(I6714A),.A1(g201A));
NAND2_X1 U_g2310A (.ZN(g2310A),.A2(g605A),.A1(g591A));
NAND2_X1 U_I7685A (.ZN(I7685A),.A2(I7683A),.A1(g3460A));
NAND2_X1 U_g3056A (.ZN(g3056A),.A2(g599A),.A1(g2374A));
NAND2_X1 U_I12108A (.ZN(I12108A),.A2(I12106A),.A1(g135A));
NAND3_X1 U_g3529A (.ZN(g3529A),.A3(g2325A),.A2(g3062A),.A1(g2310A));
NAND2_X1 U_I6747A (.ZN(I6747A),.A2(I6746A),.A1(g2938A));
NAND2_X1 U_g2236A (.ZN(g2236A),.A2(I5231A),.A1(I5230A));
NAND2_X1 U_g7584A (.ZN(g7584A),.A2(I12076A),.A1(I12075A));
NAND2_X1 U_I15870A (.ZN(I15870A),.A2(FE_OFN239_g1796A),.A1(g10291A));
NAND2_X1 U_I16067A (.ZN(I16067A),.A2(I16065A),.A1(FE_OFN237_g1806A));
NAND2_X1 U_I7562A (.ZN(I7562A),.A2(g654A),.A1(g3533A));
NAND2_X1 U_I13531A (.ZN(I13531A),.A2(I13529A),.A1(g8253A));
NAND2_X1 U_I8797A (.ZN(I8797A),.A2(I8795A),.A1(g1145A));
NAND2_X1 U_I17584A (.ZN(I17584A),.A2(g11515A),.A1(g11217A));
NAND2_X1 U_I11936A (.ZN(I11936A),.A2(I11935A),.A1(g5857A));
NAND2_X1 U_I15257A (.ZN(I15257A),.A2(I15256A),.A1(g9974A));
NAND2_X1 U_g8402A (.ZN(g8402A),.A2(I13506A),.A1(I13505A));
NAND3_X1 U_g8824A (.ZN(g8824A),.A3(g8512A),.A2(g8501A),.A1(g8502A));
NAND2_X1 U_I6186A (.ZN(I6186A),.A2(g466A),.A1(g2511A));
NAND2_X1 U_g11496A (.ZN(g11496A),.A2(I17505A),.A1(I17504A));
NAND2_X1 U_I16001A (.ZN(I16001A),.A2(I15999A),.A1(FE_OFN247_g1771A));
NAND2_X1 U_I6125A (.ZN(I6125A),.A2(I6124A),.A1(g2215A));
NAND2_X1 U_I11909A (.ZN(I11909A),.A2(I11907A),.A1(g1474A));
NAND2_X1 U_I12040A (.ZN(I12040A),.A2(I12038A),.A1(g1466A));
NAND2_X1 U_I13909A (.ZN(I13909A),.A2(I13907A),.A1(g1432A));
NAND2_X1 U_g3625A (.ZN(g3625A),.A2(I6772A),.A1(I6771A));
NAND2_X1 U_I11908A (.ZN(I11908A),.A2(I11907A),.A1(g5838A));
NAND2_X1 U_g10470A (.ZN(g10470A),.A2(I16009A),.A1(I16008A));
NAND2_X1 U_I13908A (.ZN(I13908A),.A2(I13907A),.A1(g8265A));
NAND2_X1 U_g3813A (.ZN(g3813A),.A2(I7035A),.A1(I7034A));
NAND2_X1 U_I8650A (.ZN(I8650A),.A2(g778A),.A1(g4824A));
NAND2_X1 U_g6207A (.ZN(g6207A),.A2(I9948A),.A1(I9947A));
NAND2_X1 U_I16066A (.ZN(I16066A),.A2(I16065A),.A1(g10428A));
NAND2_X1 U_g2948A (.ZN(g2948A),.A2(I6145A),.A1(I6144A));
NAND2_X1 U_I11242A (.ZN(I11242A),.A2(I11241A),.A1(g6760A));
NAND2_X1 U_g10467A (.ZN(g10467A),.A2(I15994A),.A1(I15993A));
NAND2_X1 U_I6187A (.ZN(I6187A),.A2(I6186A),.A1(g2511A));
NAND2_X1 U_g6488A (.ZN(g6488A),.A2(g6019A),.A1(g6027A));
NAND2_X1 U_I5500A (.ZN(I5500A),.A2(g1007A),.A1(g1255A));
NAND2_X1 U_I11974A (.ZN(I11974A),.A2(I11973A),.A1(g5852A));
NAND2_X1 U_I12062A (.ZN(I12062A),.A2(I12060A),.A1(g1478A));
NAND2_X1 U_g5300A (.ZN(g5300A),.A2(I8772A),.A1(I8771A));
NAND2_X1 U_I5184A (.ZN(I5184A),.A2(g1515A),.A1(g1415A));
NAND2_X1 U_I13293A (.ZN(I13293A),.A2(g8161A),.A1(g1882A));
NAND2_X1 U_I6200A (.ZN(I6200A),.A2(I6199A),.A1(g2525A));
NAND2_X1 U_I13265A (.ZN(I13265A),.A2(g8154A),.A1(g1909A));
NAND2_X1 U_I5024A (.ZN(I5024A),.A2(I5023A),.A1(g995A));
NAND2_X1 U_I7863A (.ZN(I7863A),.A2(g774A),.A1(g4099A));
NAND2_X1 U_g8705A (.ZN(g8705A),.A2(I13992A),.A1(I13991A));
NAND2_X1 U_g8471A (.ZN(g8471A),.A2(I13661A),.A1(I13660A));
NAND2_X1 U_I15256A (.ZN(I15256A),.A2(g9968A),.A1(g9974A));
NAND2_X1 U_I6145A (.ZN(I6145A),.A2(I6143A),.A1(g646A));
NAND2_X1 U_I13992A (.ZN(I13992A),.A2(I13990A),.A1(g8688A));
NAND2_X1 U_I11510A (.ZN(I11510A),.A2(I11508A),.A1(FE_OFN237_g1806A));
NAND2_X1 U_g10853A (.ZN(g10853A),.A2(g5034A),.A1(g10731A));
NAND2_X1 U_I5231A (.ZN(I5231A),.A2(I5229A),.A1(g148A));
NAND2_X1 U_I12047A (.ZN(I12047A),.A2(I12045A),.A1(g1486A));
NAND2_X1 U_I10771A (.ZN(I10771A),.A2(I10769A),.A1(g1801A));
NAND2_X1 U_g10477A (.ZN(g10477A),.A2(I16046A),.A1(I16045A));
NAND2_X1 U_g7582A (.ZN(g7582A),.A2(I12062A),.A1(I12061A));
NAND2_X1 U_I5104A (.ZN(I5104A),.A2(g435A),.A1(g431A));
NAND2_X1 U_g8409A (.ZN(g8409A),.A2(I13531A),.A1(I13530A));
NAND2_X1 U_I6447A (.ZN(I6447A),.A2(FE_OFN236_g1776A),.A1(g2264A));
NAND2_X1 U_I4956A (.ZN(I4956A),.A2(I4954A),.A1(g327A));
NAND2_X1 U_I5613A (.ZN(I5613A),.A2(I5611A),.A1(g1284A));
NAND2_X1 U_I8481A (.ZN(I8481A),.A2(I8479A),.A1(g3530A));
NAND2_X1 U_g5278A (.ZN(g5278A),.A2(I8740A),.A1(I8739A));
NAND2_X1 U_I6880A (.ZN(I6880A),.A2(I6879A),.A1(g3301A));
NAND2_X1 U_I15431A (.ZN(I15431A),.A2(I15430A),.A1(g10001A));
NAND2_X1 U_g5548A (.ZN(g5548A),.A2(FE_OFN223_g4401A),.A1(g1840A));
NAND4_X1 U_g7671A (.ZN(g7671A),.A4(FE_OFN96_g2169A),.A3(FE_OFN91_g2172A),.A2(g2175A),.A1(g2178A));
NAND2_X1 U_I12020A (.ZN(I12020A),.A2(I12019A),.A1(g6049A));
NAND2_X1 U_g10665A (.ZN(g10665A),.A2(I16332A),.A1(I16331A));
NAND2_X1 U_I16469A (.ZN(I16469A),.A2(I16467A),.A1(g10518A));
NAND2_X1 U_I5014A (.ZN(I5014A),.A2(I5013A),.A1(g1007A));
NAND2_X1 U_I13523A (.ZN(I13523A),.A2(I13521A),.A1(g8249A));
NAND2_X1 U_I16039A (.ZN(I16039A),.A2(I16037A),.A1(FE_OFN252_g1791A));
NAND2_X1 U_I16468A (.ZN(I16468A),.A2(I16467A),.A1(g10716A));
NAND2_X1 U_I12046A (.ZN(I12046A),.A2(I12045A),.A1(g5814A));
NAND2_X1 U_g4476A (.ZN(g4476A),.A2(g3071A),.A1(g3807A));
NAND2_X1 U_g10476A (.ZN(g10476A),.A2(I16039A),.A1(I16038A));
NAND2_X1 U_I16038A (.ZN(I16038A),.A2(I16037A),.A1(g10363A));
NAND2_X1 U_I8676A (.ZN(I8676A),.A2(g1027A),.A1(g4374A));
NAND2_X1 U_I12113A (.ZN(I12113A),.A2(g162A),.A1(g6002A));
NAND2_X1 U_I8761A (.ZN(I8761A),.A2(g1129A),.A1(g4616A));
NAND2_X1 U_g3204A (.ZN(g3204A),.A2(g2061A),.A1(g2571A));
NAND2_X1 U_I15993A (.ZN(I15993A),.A2(I15992A),.A1(g10430A));
NAND2_X1 U_I5036A (.ZN(I5036A),.A2(I5034A),.A1(g1019A));
NAND2_X1 U_I14263A (.ZN(I14263A),.A2(g1814A),.A1(g8843A));
NAND2_X1 U_g8298A (.ZN(g8298A),.A2(I13250A),.A1(I13249A));
NAND2_X1 U_I5135A (.ZN(I5135A),.A2(g525A),.A1(g521A));
NAND2_X1 U_g2405A (.ZN(g2405A),.A2(I5486A),.A1(I5485A));
NAND2_X1 U_I7034A (.ZN(I7034A),.A2(I7033A),.A1(g3089A));
NAND2_X1 U_I15443A (.ZN(I15443A),.A2(I15441A),.A1(g10007A));
NAND2_X1 U_I6166A (.ZN(I6166A),.A2(g153A),.A1(g2236A));
NAND2_X1 U_I8624A (.ZN(I8624A),.A2(g511A),.A1(g4267A));
NAND2_X1 U_I16015A (.ZN(I16015A),.A2(g1781A),.A1(g10441A));
NAND2_X1 U_I8677A (.ZN(I8677A),.A2(I8676A),.A1(g4374A));
NAND2_X1 U_I8576A (.ZN(I8576A),.A2(I8575A),.A1(g4234A));
NAND2_X1 U_I14613A (.ZN(I14613A),.A2(I14612A),.A1(g9204A));
NAND2_X1 U_I8716A (.ZN(I8716A),.A2(I8715A),.A1(g4601A));
NAND2_X1 U_g3530A (.ZN(g3530A),.A2(I6716A),.A1(I6715A));
NAND2_X1 U_g8405A (.ZN(g8405A),.A2(I13515A),.A1(I13514A));
NAND4_X1 U_g4104A (.ZN(g4104A),.A4(g3200A),.A3(g2439A),.A2(g3247A),.A1(g3215A));
NAND2_X1 U_I12003A (.ZN(I12003A),.A2(I12002A),.A1(g5996A));
NAND2_X1 U_g2177A (.ZN(g2177A),.A2(I5128A),.A1(I5127A));
NAND2_X1 U_g3010A (.ZN(g3010A),.A2(g2399A),.A1(g2382A));
NAND2_X1 U_g5179A (.ZN(g5179A),.A2(I8577A),.A1(I8576A));
NAND2_X1 U_I17395A (.ZN(I17395A),.A2(I17393A),.A1(g11414A));
NAND2_X1 U_g7067A (.ZN(g7067A),.A2(I11280A),.A1(I11279A));
NAND4_X1 U_g7994A (.ZN(g7994A),.A4(g7550A),.A3(FE_OFN91_g2172A),.A2(g7574A),.A1(FE_OFN88_g2178A));
NAND2_X1 U_I6167A (.ZN(I6167A),.A2(I6166A),.A1(g2236A));
NAND2_X1 U_I5265A (.ZN(I5265A),.A2(I5263A),.A1(g461A));
NAND2_X1 U_I6989A (.ZN(I6989A),.A2(I6988A),.A1(g2760A));
NAND2_X1 U_I13274A (.ZN(I13274A),.A2(I13272A),.A1(g8158A));
NAND2_X1 U_I10507A (.ZN(I10507A),.A2(g786A),.A1(g6221A));
NAND2_X1 U_I13530A (.ZN(I13530A),.A2(I13529A),.A1(g704A));
NAND2_X1 U_I5164A (.ZN(I5164A),.A2(g1499A),.A1(g1508A));
NAND2_X1 U_g9107A (.ZN(g9107A),.A2(I14444A),.A1(I14443A));
NAND2_X1 U_I9559A (.ZN(I9559A),.A2(I9557A),.A1(g782A));
NAND2_X1 U_I8577A (.ZN(I8577A),.A2(I8575A),.A1(g496A));
NAND2_X1 U_g2510A (.ZN(g2510A),.A2(I5593A),.A1(I5592A));
NAND2_X1 U_g8177A (.ZN(g8177A),.A2(I13078A),.A1(I13077A));
NAND2_X1 U_I8717A (.ZN(I8717A),.A2(I8715A),.A1(g4052A));
NAND2_X1 U_I5296A (.ZN(I5296A),.A2(I5295A),.A1(g794A));
NAND2_X1 U_g5209A (.ZN(g5209A),.A2(I8626A),.A1(I8625A));
NAND4_X1 U_g7950A (.ZN(g7950A),.A4(FE_OFN96_g2169A),.A3(g7562A),.A2(g7574A),.A1(g6941A));
NAND2_X1 U_g2088A (.ZN(g2088A),.A2(I4912A),.A1(I4911A));
NAND2_X1 U_I16000A (.ZN(I16000A),.A2(I15999A),.A1(g10432A));
NAND2_X1 U_I5371A (.ZN(I5371A),.A2(g976A),.A1(g971A));
NAND2_X1 U_g2215A (.ZN(g2215A),.A2(I5186A),.A1(I5185A));
NAND2_X1 U_g7101A (.ZN(g7101A),.A2(g2364A),.A1(g6617A));
NAND2_X1 U_I5675A (.ZN(I5675A),.A2(g1223A),.A1(g1218A));
NAND2_X1 U_I8544A (.ZN(I8544A),.A2(I8543A),.A1(g4218A));
NAND2_X1 U_g6577A (.ZN(g6577A),.A2(I10521A),.A1(I10520A));
NAND2_X1 U_I5297A (.ZN(I5297A),.A2(I5295A),.A1(g798A));
NAND2_X1 U_I13537A (.ZN(I13537A),.A2(g8157A),.A1(g658A));
NAND2_X1 U_I13283A (.ZN(I13283A),.A2(g8159A),.A1(g1927A));
NAND2_X1 U_g4749A (.ZN(g4749A),.A2(g2061A),.A1(g3710A));
NAND2_X1 U_I11982A (.ZN(I11982A),.A2(I11980A),.A1(g1482A));
NAND2_X1 U_I8514A (.ZN(I8514A),.A2(I8513A),.A1(g4873A));
NAND2_X1 U_I13091A (.ZN(I13091A),.A2(I13089A),.A1(g1840A));
NAND2_X1 U_g2943A (.ZN(g2943A),.A2(I6126A),.A1(I6125A));
NAND2_X1 U_I15908A (.ZN(I15908A),.A2(I15906A),.A1(g10302A));
NAND2_X1 U_I6879A (.ZN(I6879A),.A2(g1351A),.A1(g3301A));
NAND2_X1 U_I8763A (.ZN(I8763A),.A2(I8761A),.A1(g1129A));
NAND2_X1 U_I5449A (.ZN(I5449A),.A2(g991A),.A1(g1235A));
NAND3_X1 U_g8825A (.ZN(g8825A),.A3(g8506A),.A2(g8738A),.A1(g8502A));
NAND2_X1 U_I16007A (.ZN(I16007A),.A2(FE_OFN236_g1776A),.A1(g10434A));
NAND2_X1 U_I5865A (.ZN(I5865A),.A2(g2105A),.A1(g2107A));
NAND2_X1 U_I5604A (.ZN(I5604A),.A2(g1153A),.A1(g1149A));
NAND2_X1 U_g2433A (.ZN(g2433A),.A2(I5518A),.A1(I5517A));
NAND2_X1 U_I6111A (.ZN(I6111A),.A2(I6109A),.A1(g1494A));
NAND2_X1 U_g2096A (.ZN(g2096A),.A2(I4930A),.A1(I4929A));
NAND2_X1 U_I13522A (.ZN(I13522A),.A2(I13521A),.A1(g695A));
NAND2_X1 U_I10770A (.ZN(I10770A),.A2(I10769A),.A1(g5944A));
NAND2_X1 U_g6027A (.ZN(g6027A),.A2(FE_OFN200_g4921A),.A1(g4566A));
NAND4_X1 U_g7992A (.ZN(g7992A),.A4(FE_OFN96_g2169A),.A3(FE_OFN91_g2172A),.A2(g7574A),.A1(FE_OFN88_g2178A));
NAND2_X1 U_I5539A (.ZN(I5539A),.A2(I5538A),.A1(g1270A));
NAND2_X1 U_I17394A (.ZN(I17394A),.A2(I17393A),.A1(g11415A));
NAND2_X1 U_I13553A (.ZN(I13553A),.A2(I13552A),.A1(g668A));
NAND2_X1 U_I8642A (.ZN(I8642A),.A2(I8640A),.A1(g516A));
NAND2_X1 U_g7573A (.ZN(g7573A),.A2(I12047A),.A1(I12046A));
NAND2_X1 U_g11416A (.ZN(g11416A),.A2(I17297A),.A1(I17296A));
NAND2_X1 U_g6003A (.ZN(g6003A),.A2(g5548A),.A1(g5552A));
NAND2_X1 U_g8934A (.ZN(g8934A),.A2(I14279A),.A1(I14278A));
NAND2_X1 U_I15992A (.ZN(I15992A),.A2(g2677A),.A1(g10430A));
NAND2_X1 U_I7683A (.ZN(I7683A),.A2(g3460A),.A1(g1023A));
NAND2_X1 U_I4910A (.ZN(I4910A),.A2(g318A),.A1(g386A));
NAND4_X1 U_g3209A (.ZN(g3209A),.A4(g2571A),.A3(g2564A),.A2(g2061A),.A1(g2550A));
NAND2_X1 U_I6794A (.ZN(I6794A),.A2(I6792A),.A1(g143A));
NAND2_X1 U_I10521A (.ZN(I10521A),.A2(I10519A),.A1(g822A));
NAND2_X1 U_I5486A (.ZN(I5486A),.A2(I5484A),.A1(g1011A));
NAND2_X1 U_I15442A (.ZN(I15442A),.A2(I15441A),.A1(g10013A));
NAND2_X1 U_g6858A (.ZN(g6858A),.A2(I10932A),.A1(I10931A));
NAND2_X1 U_I5185A (.ZN(I5185A),.A2(I5184A),.A1(g1415A));
NAND2_X1 U_g5304A (.ZN(g5304A),.A2(I8780A),.A1(I8779A));
NAND2_X1 U_g2354A (.ZN(g2354A),.A2(g1520A),.A1(g1515A));
NAND2_X1 U_I15615A (.ZN(I15615A),.A2(g10153A),.A1(g10043A));
NAND2_X1 U_I17281A (.ZN(I17281A),.A2(g11219A),.A1(g11221A));
NAND2_X1 U_I5470A (.ZN(I5470A),.A2(I5468A),.A1(g999A));
NAND2_X1 U_I11509A (.ZN(I11509A),.A2(I11508A),.A1(g6580A));
NAND2_X1 U_I5025A (.ZN(I5025A),.A2(I5023A),.A1(g1275A));
NAND2_X1 U_I11508A (.ZN(I11508A),.A2(g1806A),.A1(g6580A));
NAND2_X1 U_I15430A (.ZN(I15430A),.A2(g9995A),.A1(g10001A));
NAND2_X1 U_I14612A (.ZN(I14612A),.A2(g611A),.A1(g9204A));
NAND2_X1 U_g4675A (.ZN(g4675A),.A2(g3247A),.A1(g4073A));
NAND2_X1 U_I14272A (.ZN(I14272A),.A2(I14270A),.A1(g1822A));
NAND2_X1 U_g2979A (.ZN(g2979A),.A2(I6209A),.A1(I6208A));
NAND2_X1 U_I17290A (.ZN(I17290A),.A2(I17288A),.A1(g11223A));
NAND2_X1 U_g5269A (.ZN(g5269A),.A2(I8717A),.A1(I8716A));
NAND2_X1 U_g4297A (.ZN(g4297A),.A2(I7564A),.A1(I7563A));
NAND2_X1 U_I12002A (.ZN(I12002A),.A2(g153A),.A1(g5996A));
NAND2_X1 U_I5006A (.ZN(I5006A),.A2(I5005A),.A1(g421A));
NAND2_X1 U_I12128A (.ZN(I12128A),.A2(I12126A),.A1(g170A));
NAND2_X1 U_I5105A (.ZN(I5105A),.A2(I5104A),.A1(g431A));
NAND2_X1 U_I6323A (.ZN(I6323A),.A2(I6322A),.A1(g2050A));
NAND2_X1 U_g7588A (.ZN(g7588A),.A2(I12094A),.A1(I12093A));
NAND2_X1 U_I6666A (.ZN(I6666A),.A2(I6664A),.A1(g2776A));
NAND2_X1 U_g3623A (.ZN(g3623A),.A2(I6762A),.A1(I6761A));
NAND2_X1 U_I5373A (.ZN(I5373A),.A2(I5371A),.A1(g976A));
NAND2_X1 U_I8529A (.ZN(I8529A),.A2(I8527A),.A1(g481A));
NAND2_X1 U_I5283A (.ZN(I5283A),.A2(I5282A),.A1(g758A));
NAND2_X1 U_I7224A (.ZN(I7224A),.A2(I7223A),.A1(g2981A));
NAND2_X1 U_I5007A (.ZN(I5007A),.A2(I5005A),.A1(g312A));
NAND2_X1 U_I5459A (.ZN(I5459A),.A2(g1003A),.A1(g1240A));
NAND2_X1 U_I17297A (.ZN(I17297A),.A2(I17295A),.A1(g11227A));
NAND3_X1 U_g8746A (.ZN(g8746A),.A3(g46A),.A2(g47A),.A1(g8617A));
NAND2_X1 U_I6143A (.ZN(I6143A),.A2(g646A),.A1(g1976A));
NAND2_X1 U_I5015A (.ZN(I5015A),.A2(I5013A),.A1(g1011A));
NAND2_X1 U_g8932A (.ZN(g8932A),.A2(I14265A),.A1(I14264A));
NAND2_X1 U_I16073A (.ZN(I16073A),.A2(I16072A),.A1(g845A));
NAND2_X1 U_I6988A (.ZN(I6988A),.A2(g986A),.A1(g2760A));
NAND2_X1 U_g3205A (.ZN(g3205A),.A2(g2571A),.A1(g1814A));
NAND2_X1 U_I8652A (.ZN(I8652A),.A2(I8650A),.A1(g778A));
NAND2_X1 U_I9558A (.ZN(I9558A),.A2(I9557A),.A1(g5598A));
NAND2_X1 U_I5203A (.ZN(I5203A),.A2(I5202A),.A1(g369A));
NAND2_X1 U_g7533A (.ZN(g7533A),.A2(I11937A),.A1(I11936A));
NAND2_X1 U_g3634A (.ZN(g3634A),.A2(I6807A),.A1(I6806A));
NAND2_X1 U_I6792A (.ZN(I6792A),.A2(g143A),.A1(g2959A));
NAND2_X1 U_g3304A (.ZN(g3304A),.A2(I6469A),.A1(I6468A));
NAND2_X1 U_I12145A (.ZN(I12145A),.A2(I12143A),.A1(g158A));
NAND2_X1 U_g7596A (.ZN(g7596A),.A2(I12128A),.A1(I12127A));
NAND2_X1 U_I13302A (.ZN(I13302A),.A2(I13300A),.A1(g8162A));
NAND2_X1 U_I5502A (.ZN(I5502A),.A2(I5500A),.A1(g1007A));
NAND2_X1 U_I9574A (.ZN(I9574A),.A2(g818A),.A1(g5608A));
NAND2_X1 U_g3273A (.ZN(g3273A),.A2(I6449A),.A1(I6448A));
NAND2_X1 U_I8670A (.ZN(I8670A),.A2(I8669A),.A1(g4831A));
NAND2_X1 U_I7035A (.ZN(I7035A),.A2(I7033A),.A1(g1868A));
NAND2_X1 U_I15453A (.ZN(I15453A),.A2(I15451A),.A1(g10019A));
NAND2_X1 U_I8625A (.ZN(I8625A),.A2(I8624A),.A1(g4267A));
NAND2_X1 U_I7876A (.ZN(I7876A),.A2(I7875A),.A1(g4109A));
NAND2_X1 U_I14203A (.ZN(I14203A),.A2(I14202A),.A1(g8825A));
NAND2_X1 U_I15607A (.ZN(I15607A),.A2(g10144A),.A1(g10149A));
NAND2_X1 U_g2274A (.ZN(g2274A),.A2(I5325A),.A1(I5324A));
NAND2_X1 U_I8740A (.ZN(I8740A),.A2(I8738A),.A1(g1121A));
NAND2_X1 U_I17296A (.ZN(I17296A),.A2(I17295A),.A1(g11229A));
NAND2_X1 U_g10507A (.ZN(g10507A),.A2(g5859A),.A1(g10434A));
NAND2_X1 U_g2325A (.ZN(g2325A),.A2(g617A),.A1(g611A));
NAND2_X1 U_I8606A (.ZN(I8606A),.A2(I8604A),.A1(g506A));
NAND2_X1 U_I12087A (.ZN(I12087A),.A2(I12085A),.A1(g1470A));
NAND2_X1 U_I13249A (.ZN(I13249A),.A2(I13248A),.A1(g1891A));
NAND2_X1 U_I13248A (.ZN(I13248A),.A2(g8148A),.A1(g1891A));
NAND2_X1 U_I13552A (.ZN(I13552A),.A2(g8262A),.A1(g668A));
NAND2_X1 U_g2106A (.ZN(g2106A),.A2(I4980A),.A1(I4979A));
NAND2_X1 U_I12069A (.ZN(I12069A),.A2(I12067A),.A1(g139A));
NAND2_X1 U_g9204A (.ZN(g9204A),.A2(g8942A),.A1(g6019A));
NAND2_X1 U_I12068A (.ZN(I12068A),.A2(I12067A),.A1(g6045A));
NAND2_X1 U_I17503A (.ZN(I17503A),.A2(g5269A),.A1(g11430A));
NAND2_X1 U_I7877A (.ZN(I7877A),.A2(I7875A),.A1(g810A));
NAND2_X1 U_I5165A (.ZN(I5165A),.A2(I5164A),.A1(g1508A));
NAND2_X1 U_g6740A (.ZN(g6740A),.A2(g2550A),.A1(g6131A));
NAND2_X1 U_I6289A (.ZN(I6289A),.A2(I6287A),.A1(g981A));
NAND2_X1 U_I6777A (.ZN(I6777A),.A2(g650A),.A1(g2892A));
NAND2_X1 U_g5171A (.ZN(g5171A),.A2(I8563A),.A1(I8562A));
NAND2_X1 U_I15891A (.ZN(I15891A),.A2(I15890A),.A1(g853A));
NAND2_X1 U_I13090A (.ZN(I13090A),.A2(I13089A),.A1(g8006A));
NAND2_X1 U_g11474A (.ZN(g11474A),.A2(I17461A),.A1(I17460A));
NAND4_X1 U_g7942A (.ZN(g7942A),.A4(g7550A),.A3(g7562A),.A2(FE_OFN80_g2175A),.A1(g6941A));
NAND2_X1 U_I5538A (.ZN(I5538A),.A2(g1023A),.A1(g1270A));
NAND2_X1 U_I7563A (.ZN(I7563A),.A2(I7562A),.A1(g3533A));
NAND2_X1 U_I13513A (.ZN(I13513A),.A2(g8248A),.A1(g686A));
NAND2_X1 U_g2107A (.ZN(g2107A),.A2(I4987A),.A1(I4986A));
NAND2_X1 U_g2223A (.ZN(g2223A),.A2(I5204A),.A1(I5203A));
NAND2_X1 U_I13505A (.ZN(I13505A),.A2(I13504A),.A1(g677A));
NAND2_X1 U_I6209A (.ZN(I6209A),.A2(I6207A),.A1(g802A));
NAND2_X1 U_I12086A (.ZN(I12086A),.A2(I12085A),.A1(g5842A));
NAND2_X1 U_I8545A (.ZN(I8545A),.A2(I8543A),.A1(g486A));
NAND2_X1 U_I8180A (.ZN(I8180A),.A2(I8178A),.A1(FE_OFN253_g1786A));
NAND2_X1 U_g2115A (.ZN(g2115A),.A2(I5015A),.A1(I5014A));
NAND2_X1 U_I8591A (.ZN(I8591A),.A2(I8589A),.A1(g501A));
NAND2_X1 U_I10931A (.ZN(I10931A),.A2(I10930A),.A1(g5863A));
NAND2_X1 U_I17402A (.ZN(I17402A),.A2(I17400A),.A1(g11416A));
NAND2_X1 U_g8307A (.ZN(g8307A),.A2(I13295A),.A1(I13294A));
NAND2_X1 U_I12144A (.ZN(I12144A),.A2(I12143A),.A1(g6000A));
NAND2_X1 U_I10520A (.ZN(I10520A),.A2(I10519A),.A1(g6231A));
NAND2_X1 U_I5263A (.ZN(I5263A),.A2(FE_OFN254_g461A),.A1(g456A));
NAND2_X1 U_g8757A (.ZN(g8757A),.A2(FE_OFN223_g4401A),.A1(g8599A));
NAND2_X1 U_I6714A (.ZN(I6714A),.A2(g201A),.A1(g2961A));
NAND2_X1 U_I14211A (.ZN(I14211A),.A2(I14209A),.A1(g599A));
NAND2_X1 U_I8515A (.ZN(I8515A),.A2(I8513A),.A1(g3513A));
NAND2_X1 U_g2272A (.ZN(g2272A),.A2(I5317A),.A1(I5316A));
NAND2_X1 U_I9946A (.ZN(I9946A),.A2(g1796A),.A1(g5233A));
NAND2_X1 U_I8750A (.ZN(I8750A),.A2(g1125A),.A1(g4613A));
NAND2_X1 U_I5605A (.ZN(I5605A),.A2(I5604A),.A1(g1149A));
NAND2_X1 U_g8880A (.ZN(g8880A),.A2(I14204A),.A1(I14203A));
NAND2_X1 U_I16051A (.ZN(I16051A),.A2(g10434A),.A1(g837A));
NAND2_X1 U_I16072A (.ZN(I16072A),.A2(g10438A),.A1(g845A));
NAND2_X1 U_g10440A (.ZN(g10440A),.A2(g6037A),.A1(g10360A));
NAND2_X1 U_g8612A (.ZN(g8612A),.A2(I13859A),.A1(I13858A));
NAND2_X1 U_I15872A (.ZN(I15872A),.A2(I15870A),.A1(FE_OFN239_g1796A));
NAND2_X1 U_I8528A (.ZN(I8528A),.A2(I8527A),.A1(g4879A));
NAND2_X1 U_g8629A (.ZN(g8629A),.A2(I13902A),.A1(I13901A));
NAND4_X1 U_g8542A (.ZN(g8542A),.A4(g8390A),.A3(g1814A),.A2(g1828A),.A1(g2571A));
NAND2_X1 U_I9947A (.ZN(I9947A),.A2(I9946A),.A1(g5233A));
NAND2_X1 U_I6838A (.ZN(I6838A),.A2(I6836A),.A1(g806A));
NAND2_X1 U_g7583A (.ZN(g7583A),.A2(I12069A),.A1(I12068A));
NAND2_X1 U_g4803A (.ZN(g4803A),.A2(FE_OFN325_g18A),.A1(g3664A));
NAND2_X1 U_I17307A (.ZN(I17307A),.A2(I17305A),.A1(g11231A));
NAND2_X1 U_g4538A (.ZN(g4538A),.A2(g2399A),.A1(g3475A));
NAND2_X1 U_I15452A (.ZN(I15452A),.A2(I15451A),.A1(g10025A));
NAND2_X1 U_I13857A (.ZN(I13857A),.A2(g1448A),.A1(g8270A));
NAND2_X1 U_I14202A (.ZN(I14202A),.A2(g591A),.A1(g8825A));
NAND2_X1 U_I13765A (.ZN(I13765A),.A2(g8417A),.A1(g731A));
NAND2_X1 U_g2260A (.ZN(g2260A),.A2(I5297A),.A1(I5296A));
NAND4_X1 U_g7986A (.ZN(g7986A),.A4(g7550A),.A3(g2172A),.A2(FE_OFN80_g2175A),.A1(FE_OFN88_g2178A));
NAND2_X1 U_g5226A (.ZN(g5226A),.A2(I8671A),.A1(I8670A));
NAND2_X1 U_g8512A (.ZN(g8512A),.A2(g8366A),.A1(g3723A));
NAND2_X1 U_I16046A (.ZN(I16046A),.A2(I16044A),.A1(g10432A));
NAND2_X1 U_I13504A (.ZN(I13504A),.A2(g8247A),.A1(g677A));
NAND2_X1 U_g10447A (.ZN(g10447A),.A2(g5360A),.A1(g10363A));
NAND2_X1 U_g2167A (.ZN(g2167A),.A2(I5106A),.A1(I5105A));
NAND2_X1 U_I8804A (.ZN(I8804A),.A2(I8803A),.A1(g4677A));
NAND2_X1 U_g10472A (.ZN(g10472A),.A2(I16017A),.A1(I16016A));
NAND2_X1 U_I17487A (.ZN(I17487A),.A2(I17485A),.A1(g11474A));
NAND2_X1 U_I4995A (.ZN(I4995A),.A2(g309A),.A1(g416A));
NAND2_X1 U_I12093A (.ZN(I12093A),.A2(I12092A),.A1(g5810A));
NAND4_X1 U_g7987A (.ZN(g7987A),.A4(FE_OFN96_g2169A),.A3(g7562A),.A2(FE_OFN80_g2175A),.A1(FE_OFN88_g2178A));
NAND2_X1 U_g5227A (.ZN(g5227A),.A2(I8678A),.A1(I8677A));
NAND2_X1 U_I5126A (.ZN(I5126A),.A2(g1389A),.A1(g1386A));
NAND2_X1 U_g2321A (.ZN(g2321A),.A2(I5373A),.A1(I5372A));
NAND2_X1 U_g7547A (.ZN(g7547A),.A2(I11975A),.A1(I11974A));
NAND2_X1 U_I17306A (.ZN(I17306A),.A2(I17305A),.A1(g11232A));
NAND3_X1 U_g6548A (.ZN(g6548A),.A3(g6122A),.A2(g6124A),.A1(g826A));
NAND2_X1 U_I11995A (.ZN(I11995A),.A2(g127A),.A1(g6035A));
NAND2_X1 U_I7225A (.ZN(I7225A),.A2(I7223A),.A1(g1781A));
NAND2_X1 U_I11261A (.ZN(I11261A),.A2(g826A),.A1(g6775A));
NAND3_X1 U_g8843A (.ZN(g8843A),.A3(g8545A),.A2(g8757A),.A1(g8542A));
NAND2_X1 U_g2938A (.ZN(g2938A),.A2(I6111A),.A1(I6110A));
NAND2_X1 U_I4942A (.ZN(I4942A),.A2(I4941A),.A1(g396A));
NAND2_X1 U_g10394A (.ZN(g10394A),.A2(I15900A),.A1(I15899A));
NAND2_X1 U_g8549A (.ZN(g8549A),.A2(g8390A),.A1(g5527A));
NAND2_X1 U_g3070A (.ZN(g3070A),.A2(g1206A),.A1(g2016A));
NAND2_X1 U_I4954A (.ZN(I4954A),.A2(g327A),.A1(g401A));
NAND2_X1 U_I5023A (.ZN(I5023A),.A2(g1275A),.A1(g995A));
NAND2_X1 U_g10446A (.ZN(g10446A),.A2(g5350A),.A1(g10438A));
NAND2_X1 U_I16081A (.ZN(I16081A),.A2(I16079A),.A1(g10363A));
NAND2_X1 U_I8641A (.ZN(I8641A),.A2(I8640A),.A1(g4278A));
NAND2_X1 U_I6178A (.ZN(I6178A),.A2(I6176A),.A1(g197A));
NAND2_X1 U_I12075A (.ZN(I12075A),.A2(I12074A),.A1(g6015A));
NAND2_X1 U_I5127A (.ZN(I5127A),.A2(I5126A),.A1(g1386A));
NAND2_X1 U_I5451A (.ZN(I5451A),.A2(I5449A),.A1(g991A));
NAND2_X1 U_g4168A (.ZN(g4168A),.A2(I7323A),.A1(I7322A));
NAND2_X1 U_I6288A (.ZN(I6288A),.A2(I6287A),.A1(g2091A));
NAND2_X1 U_I8179A (.ZN(I8179A),.A2(I8178A),.A1(g3685A));
NAND2_X1 U_I4912A (.ZN(I4912A),.A2(I4910A),.A1(g318A));
NAND2_X1 U_I6805A (.ZN(I6805A),.A2(g471A),.A1(g3268A));
NAND3_X1 U_g3766A (.ZN(g3766A),.A3(g2493A),.A2(g3222A),.A1(g2439A));
NAND2_X1 U_g3087A (.ZN(g3087A),.A2(I6289A),.A1(I6288A));
NAND2_X1 U_I17486A (.ZN(I17486A),.A2(I17485A),.A1(g11233A));
NAND2_X1 U_I4929A (.ZN(I4929A),.A2(I4928A),.A1(g391A));
NAND2_X1 U_I15890A (.ZN(I15890A),.A2(g10285A),.A1(g853A));
NAND2_X1 U_I16331A (.ZN(I16331A),.A2(I16330A),.A1(g10387A));
NAND2_X1 U_I9575A (.ZN(I9575A),.A2(I9574A),.A1(g5608A));
NAND2_X1 U_I13887A (.ZN(I13887A),.A2(I13886A),.A1(g8267A));
NAND2_X1 U_g5308A (.ZN(g5308A),.A2(I8788A),.A1(I8787A));
NAND2_X1 U_I13529A (.ZN(I13529A),.A2(g8253A),.A1(g704A));
NAND2_X1 U_I6208A (.ZN(I6208A),.A2(I6207A),.A1(g5188A));
NAND2_X1 U_g5217A (.ZN(g5217A),.A2(I8642A),.A1(I8641A));
NAND2_X1 U_I5316A (.ZN(I5316A),.A2(I5315A),.A1(g1032A));
NAND2_X1 U_g2111A (.ZN(g2111A),.A2(I5007A),.A1(I5006A));
NAND2_X1 U_g10366A (.ZN(g10366A),.A2(g5392A),.A1(g10285A));
NAND2_X1 U_I5034A (.ZN(I5034A),.A2(g1019A),.A1(g1015A));
NAND2_X1 U_I13869A (.ZN(I13869A),.A2(I13867A),.A1(g1403A));
NAND2_X1 U_I13868A (.ZN(I13868A),.A2(I13867A),.A1(g8264A));
NAND2_X1 U_I15999A (.ZN(I15999A),.A2(FE_OFN247_g1771A),.A1(g10432A));
NAND2_X1 U_I13259A (.ZN(I13259A),.A2(I13258A),.A1(g1900A));
NAND4_X1 U_g3261A (.ZN(g3261A),.A4(g2202A),.A3(g2211A),.A2(g2222A),.A1(g2229A));
NAND2_X1 U_g10481A (.ZN(g10481A),.A2(I16074A),.A1(I16073A));
NAND2_X1 U_g2180A (.ZN(g2180A),.A2(I5137A),.A1(I5136A));
NAND3_X1 U_g4976A (.ZN(g4976A),.A3(g3807A),.A2(g4604A),.A1(g2310A));
NAND2_X1 U_g8506A (.ZN(g8506A),.A2(g8366A),.A1(g3475A));
NAND2_X1 U_g2380A (.ZN(g2380A),.A2(I5461A),.A1(I5460A));
NAND2_X1 U_I13258A (.ZN(I13258A),.A2(g8153A),.A1(g1900A));
NAND2_X1 U_I5013A (.ZN(I5013A),.A2(g1011A),.A1(g1007A));
NAND2_X1 U_g5196A (.ZN(g5196A),.A2(I8606A),.A1(I8605A));
NAND2_X1 U_I10930A (.ZN(I10930A),.A2(g5555A),.A1(g5863A));
NAND2_X1 U_I6770A (.ZN(I6770A),.A2(g382A),.A1(g3257A));
NAND2_X1 U_g11449A (.ZN(g11449A),.A2(I17402A),.A1(I17401A));
NAND2_X1 U_g11448A (.ZN(g11448A),.A2(I17395A),.A1(I17394A));
NAND2_X1 U_I15717A (.ZN(I15717A),.A2(I15716A),.A1(g10231A));
NAND2_X1 U_I5317A (.ZN(I5317A),.A2(I5315A),.A1(g1027A));
NAND2_X1 U_I14210A (.ZN(I14210A),.A2(I14209A),.A1(g8824A));
NAND2_X1 U_I17569A (.ZN(I17569A),.A2(I17567A),.A1(g1610A));
NAND2_X1 U_I13878A (.ZN(I13878A),.A2(I13876A),.A1(g1444A));
NAND2_X1 U_g8545A (.ZN(g8545A),.A2(g8390A),.A1(g3710A));
NAND2_X1 U_g2515A (.ZN(g2515A),.A2(I5606A),.A1(I5605A));
NAND2_X1 U_I14443A (.ZN(I14443A),.A2(I14442A),.A1(g8970A));
NAND2_X1 U_g7557A (.ZN(g7557A),.A2(I11997A),.A1(I11996A));
NAND2_X1 U_g8180A (.ZN(g8180A),.A2(I13091A),.A1(I13090A));
NAND2_X1 U_I14279A (.ZN(I14279A),.A2(I14277A),.A1(g1828A));
NAND2_X1 U_I17568A (.ZN(I17568A),.A2(I17567A),.A1(g11496A));
NAND2_X1 U_I13886A (.ZN(I13886A),.A2(g1440A),.A1(g8267A));
NAND2_X1 U_I7322A (.ZN(I7322A),.A2(I7321A),.A1(g3047A));
NAND2_X1 U_I6990A (.ZN(I6990A),.A2(I6988A),.A1(g986A));
NAND2_X1 U_I14278A (.ZN(I14278A),.A2(I14277A),.A1(g8847A));
NAND2_X1 U_I7033A (.ZN(I7033A),.A2(g1868A),.A1(g3089A));
NAND2_X1 U_I9006A (.ZN(I9006A),.A2(FE_OFN252_g1791A),.A1(g4492A));
NAND2_X1 U_g8507A (.ZN(g8507A),.A2(g8366A),.A1(g3738A));
NAND2_X1 U_I5460A (.ZN(I5460A),.A2(I5459A),.A1(g1240A));
NAND2_X1 U_g4588A (.ZN(g4588A),.A2(FE_OFN325_g18A),.A1(g3440A));
NAND2_X1 U_I4986A (.ZN(I4986A),.A2(I4985A),.A1(g999A));
NAND3_X1 U_g3247A (.ZN(g3247A),.A3(g2571A),.A2(g2564A),.A1(g1828A));
NAND2_X1 U_I8651A (.ZN(I8651A),.A2(I8650A),.A1(g4824A));
NAND2_X1 U_I13545A (.ZN(I13545A),.A2(I13544A),.A1(g713A));
NAND2_X1 U_g8628A (.ZN(g8628A),.A2(I13895A),.A1(I13894A));
NAND2_X1 U_I6138A (.ZN(I6138A),.A2(I6136A),.A1(g378A));
NAND2_X1 U_I12074A (.ZN(I12074A),.A2(g174A),.A1(g6015A));
NAND2_X1 U_g8630A (.ZN(g8630A),.A2(I13909A),.A1(I13908A));
NAND2_X1 U_I13078A (.ZN(I13078A),.A2(I13076A),.A1(g7963A));
NAND2_X1 U_I6109A (.ZN(I6109A),.A2(g1494A),.A1(g2205A));
NAND2_X1 U_g8300A (.ZN(g8300A),.A2(I13260A),.A1(I13259A));
NAND2_X1 U_I5501A (.ZN(I5501A),.A2(I5500A),.A1(g1255A));
NAND2_X1 U_I17586A (.ZN(I17586A),.A2(I17584A),.A1(g11515A));
NAND2_X1 U_I12092A (.ZN(I12092A),.A2(g1490A),.A1(g5810A));
NAND2_X1 U_I13901A (.ZN(I13901A),.A2(I13900A),.A1(g8261A));
NAND2_X1 U_I8795A (.ZN(I8795A),.A2(g1145A),.A1(g4672A));
NAND2_X1 U_I6201A (.ZN(I6201A),.A2(I6199A),.A1(g766A));
NAND2_X1 U_I14217A (.ZN(I14217A),.A2(I14216A),.A1(g8826A));
NAND2_X1 U_I9007A (.ZN(I9007A),.A2(I9006A),.A1(g4492A));
NAND2_X1 U_I13561A (.ZN(I13561A),.A2(I13559A),.A1(g8263A));
NAND2_X1 U_I15716A (.ZN(I15716A),.A2(g10229A),.A1(g10231A));
NAND2_X1 U_I6449A (.ZN(I6449A),.A2(I6447A),.A1(FE_OFN236_g1776A));
NAND2_X1 U_I13295A (.ZN(I13295A),.A2(I13293A),.A1(g8161A));
NAND2_X1 U_I4987A (.ZN(I4987A),.A2(I4985A),.A1(g1003A));
NAND2_X1 U_I6715A (.ZN(I6715A),.A2(I6714A),.A1(g2961A));
NAND2_X1 U_I17493A (.ZN(I17493A),.A2(I17492A),.A1(g11430A));
NAND2_X1 U_I12215A (.ZN(I12215A),.A2(I12214A),.A1(g7061A));
NAND2_X1 U_g2372A (.ZN(g2372A),.A2(I5451A),.A1(I5450A));
NAND2_X1 U_g7062A (.ZN(g7062A),.A2(I11263A),.A1(I11262A));
NAND2_X1 U_g2988A (.ZN(g2988A),.A2(I6226A),.A1(I6225A));
NAND2_X1 U_I13309A (.ZN(I13309A),.A2(I13307A),.A1(g617A));
NAND2_X1 U_g8839A (.ZN(g8839A),.A2(FE_OFN223_g4401A),.A1(g8603A));
NAND2_X1 U_g2555A (.ZN(g2555A),.A2(I5677A),.A1(I5676A));
NAND2_X1 U_g3662A (.ZN(g3662A),.A2(I6827A),.A1(I6826A));
NAND2_X1 U_I13308A (.ZN(I13308A),.A2(I13307A),.A1(g8190A));
NAND2_X1 U_g2792A (.ZN(g2792A),.A2(I5880A),.A1(I5879A));
NAND2_X1 U_g4117A (.ZN(g4117A),.A2(g3061A),.A1(g3041A));
NAND2_X1 U_I8543A (.ZN(I8543A),.A2(g486A),.A1(g4218A));
NAND2_X1 U_g11549A (.ZN(g11549A),.A2(I17586A),.A1(I17585A));
NAND2_X1 U_I6881A (.ZN(I6881A),.A2(I6879A),.A1(g1351A));
NAND2_X1 U_I12138A (.ZN(I12138A),.A2(I12136A),.A1(g131A));
NAND2_X1 U_I8729A (.ZN(I8729A),.A2(I8728A),.A1(g4605A));
NAND2_X1 U_I14216A (.ZN(I14216A),.A2(g605A),.A1(g8826A));
NAND2_X1 U_g10384A (.ZN(g10384A),.A2(I15872A),.A1(I15871A));
NAND2_X1 U_I13260A (.ZN(I13260A),.A2(I13258A),.A1(g8153A));
NAND2_X1 U_g2776A (.ZN(g2776A),.A2(I5867A),.A1(I5866A));
NAND2_X1 U_I8513A (.ZN(I8513A),.A2(g3513A),.A1(g4873A));
NAND2_X1 U_I13559A (.ZN(I13559A),.A2(g8263A),.A1(g722A));
NAND2_X1 U_I8178A (.ZN(I8178A),.A2(FE_OFN253_g1786A),.A1(g3685A));
NAND2_X1 U_g3631A (.ZN(g3631A),.A2(I6794A),.A1(I6793A));
NAND2_X1 U_I6487A (.ZN(I6487A),.A2(g1227A),.A1(g2306A));
NAND2_X1 U_I16080A (.ZN(I16080A),.A2(I16079A),.A1(g849A));
NAND2_X1 U_I13893A (.ZN(I13893A),.A2(g1436A),.A1(g8266A));
NAND2_X1 U_I12115A (.ZN(I12115A),.A2(I12113A),.A1(g162A));
NAND2_X1 U_I6748A (.ZN(I6748A),.A2(I6746A),.A1(g1453A));
NAND2_X1 U_I13544A (.ZN(I13544A),.A2(g8259A),.A1(g713A));
NAND2_X1 U_I5484A (.ZN(I5484A),.A2(g1011A),.A1(g1250A));
NAND2_X1 U_I4928A (.ZN(I4928A),.A2(g321A),.A1(g391A));
NAND2_X1 U_I6226A (.ZN(I6226A),.A2(I6224A),.A1(g1346A));
NAND2_X1 U_I8805A (.ZN(I8805A),.A2(I8803A),.A1(g1113A));
NAND2_X1 U_I4930A (.ZN(I4930A),.A2(I4928A),.A1(g321A));
NAND2_X1 U_I15880A (.ZN(I15880A),.A2(I15878A),.A1(FE_OFN251_g1801A));
NAND2_X1 U_I14265A (.ZN(I14265A),.A2(I14263A),.A1(g1814A));
NAND2_X1 U_I16031A (.ZN(I16031A),.A2(I16030A),.A1(g829A));
NAND2_X1 U_g3585A (.ZN(g3585A),.A2(I6748A),.A1(I6747A));
NAND4_X1 U_g3041A (.ZN(g3041A),.A4(g2382A),.A3(g2374A),.A2(g2399A),.A1(g2364A));
NAND2_X1 U_g8933A (.ZN(g8933A),.A2(I14272A),.A1(I14271A));
NAND2_X1 U_I16330A (.ZN(I16330A),.A2(g4997A),.A1(g10387A));
NAND2_X1 U_I13267A (.ZN(I13267A),.A2(I13265A),.A1(g8154A));
NAND2_X1 U_I13294A (.ZN(I13294A),.A2(I13293A),.A1(g1882A));
NAND2_X1 U_g10231A (.ZN(g10231A),.A2(I15617A),.A1(I15616A));
NAND2_X1 U_I14442A (.ZN(I14442A),.A2(g1834A),.A1(g8970A));
NAND2_X1 U_I6793A (.ZN(I6793A),.A2(I6792A),.A1(g2959A));
NAND2_X1 U_I4966A (.ZN(I4966A),.A2(I4964A),.A1(g330A));
NAND2_X1 U_I8752A (.ZN(I8752A),.A2(I8750A),.A1(g1125A));
NAND2_X1 U_I15432A (.ZN(I15432A),.A2(I15430A),.A1(g9995A));
NAND2_X1 U_I12214A (.ZN(I12214A),.A2(g2518A),.A1(g7061A));
NAND2_X1 U_g10511A (.ZN(g10511A),.A2(g6032A),.A1(g10438A));
NAND2_X1 U_g3011A (.ZN(g3011A),.A2(g2382A),.A1(g591A));
NAND2_X1 U_g5103A (.ZN(g5103A),.A2(I8481A),.A1(I8480A));
NAND2_X1 U_I16087A (.ZN(I16087A),.A2(I16086A),.A1(g861A));
NAND2_X1 U_g3734A (.ZN(g3734A),.A2(g599A),.A1(g3039A));
NAND2_X1 U_I6664A (.ZN(I6664A),.A2(g2776A),.A1(g2792A));
NAND2_X1 U_g8882A (.ZN(g8882A),.A2(I14218A),.A1(I14217A));
NAND2_X1 U_I4955A (.ZN(I4955A),.A2(I4954A),.A1(g401A));
NAND2_X1 U_I8786A (.ZN(I8786A),.A2(g1141A),.A1(g4639A));
NAND3_X1 U_g3992A (.ZN(g3992A),.A3(g2990A),.A2(g2550A),.A1(g2571A));
NAND2_X1 U_g10480A (.ZN(g10480A),.A2(I16067A),.A1(I16066A));
NAND2_X1 U_I11915A (.ZN(I11915A),.A2(I11914A),.A1(g5803A));
NAND2_X1 U_I8770A (.ZN(I8770A),.A2(g1133A),.A1(g4619A));
NAND2_X1 U_I5516A (.ZN(I5516A),.A2(g1019A),.A1(g1260A));
NAND2_X1 U_g8541A (.ZN(g8541A),.A2(g8390A),.A1(g4001A));
NAND2_X1 U_I6188A (.ZN(I6188A),.A2(I6186A),.A1(g466A));
NAND2_X1 U_g5147A (.ZN(g5147A),.A2(I8545A),.A1(I8544A));
NAND3_X1 U_g8744A (.ZN(g8744A),.A3(I9273A),.A2(g46A),.A1(g8617A));
NAND2_X1 U_I5892A (.ZN(I5892A),.A2(I5891A),.A1(g750A));
NAND2_X1 U_g8558A (.ZN(g8558A),.A2(I13767A),.A1(I13766A));
NAND2_X1 U_I15258A (.ZN(I15258A),.A2(I15256A),.A1(g9968A));
NAND2_X1 U_I13266A (.ZN(I13266A),.A2(I13265A),.A1(g1909A));
NAND2_X1 U_I8787A (.ZN(I8787A),.A2(I8786A),.A1(g4639A));
NAND2_X1 U_I6826A (.ZN(I6826A),.A2(I6825A),.A1(g3281A));
NAND2_X1 U_I17283A (.ZN(I17283A),.A2(I17281A),.A1(g11219A));
NAND3_X1 U_g5013A (.ZN(g5013A),.A3(g3205A),.A2(g3247A),.A1(g4749A));
NAND2_X1 U_I17492A (.ZN(I17492A),.A2(g3623A),.A1(g11430A));
NAND2_X1 U_g8511A (.ZN(g8511A),.A2(g8366A),.A1(g5277A));
NAND2_X1 U_I16079A (.ZN(I16079A),.A2(g10363A),.A1(g849A));
NAND2_X1 U_I5035A (.ZN(I5035A),.A2(I5034A),.A1(g1015A));
NAND2_X1 U_I5517A (.ZN(I5517A),.A2(I5516A),.A1(g1260A));
NAND2_X1 U_I7223A (.ZN(I7223A),.A2(g1781A),.A1(g2981A));
NAND2_X1 U_I16086A (.ZN(I16086A),.A2(g10430A),.A1(g861A));
NAND2_X1 U_g5317A (.ZN(g5317A),.A2(I8797A),.A1(I8796A));
NAND2_X1 U_I15879A (.ZN(I15879A),.A2(I15878A),.A1(g10359A));
NAND2_X1 U_I15878A (.ZN(I15878A),.A2(FE_OFN251_g1801A),.A1(g10359A));
NAND2_X1 U_I12114A (.ZN(I12114A),.A2(I12113A),.A1(g6002A));
NAND2_X1 U_I12107A (.ZN(I12107A),.A2(I12106A),.A1(g6042A));
NAND2_X1 U_g2500A (.ZN(g2500A),.A2(g182A),.A1(g178A));
NAND2_X1 U_I15994A (.ZN(I15994A),.A2(I15992A),.A1(g2677A));
NAND4_X1 U_g7934A (.ZN(g7934A),.A4(g7550A),.A3(FE_OFN91_g2172A),.A2(FE_OFN80_g2175A),.A1(g6941A));
NAND2_X1 U_g10469A (.ZN(g10469A),.A2(g5999A),.A1(g10430A));
NAND2_X1 U_I14264A (.ZN(I14264A),.A2(I14263A),.A1(g8843A));
NAND2_X1 U_I6448A (.ZN(I6448A),.A2(I6447A),.A1(g2264A));
NAND2_X1 U_I13285A (.ZN(I13285A),.A2(I13283A),.A1(g8159A));
NAND2_X1 U_g10468A (.ZN(g10468A),.A2(I16001A),.A1(I16000A));
NAND2_X1 U_I6827A (.ZN(I6827A),.A2(I6825A),.A1(g770A));
NAND2_X1 U_g8623A (.ZN(g8623A),.A2(I13878A),.A1(I13877A));
NAND2_X1 U_I13900A (.ZN(I13900A),.A2(g1428A),.A1(g8261A));
NAND2_X1 U_g2795A (.ZN(g2795A),.A2(I5893A),.A1(I5892A));
NAND2_X1 U_I8575A (.ZN(I8575A),.A2(g496A),.A1(g4234A));
NAND2_X1 U_I14209A (.ZN(I14209A),.A2(g599A),.A1(g8824A));
NAND2_X1 U_I13560A (.ZN(I13560A),.A2(I13559A),.A1(g722A));
NAND2_X1 U_I8715A (.ZN(I8715A),.A2(g4052A),.A1(g4601A));
NAND2_X1 U_I8604A (.ZN(I8604A),.A2(g506A),.A1(g4259A));
NAND2_X1 U_I16017A (.ZN(I16017A),.A2(I16015A),.A1(g1781A));
NAND2_X1 U_I4941A (.ZN(I4941A),.A2(g324A),.A1(g396A));
NAND2_X1 U_g2205A (.ZN(g2205A),.A2(I5166A),.A1(I5165A));
NAND3_X1 U_g3753A (.ZN(g3753A),.A3(g2800A),.A2(g2364A),.A1(g2382A));
NAND2_X1 U_I6467A (.ZN(I6467A),.A2(g2479A),.A1(g23A));
NAND2_X1 U_I14614A (.ZN(I14614A),.A2(I14612A),.A1(g611A));
NAND2_X1 U_g2104A (.ZN(g2104A),.A2(I4966A),.A1(I4965A));
NAND2_X1 U_g2099A (.ZN(g2099A),.A2(I4943A),.A1(I4942A));
NAND2_X1 U_I16023A (.ZN(I16023A),.A2(FE_OFN253_g1786A),.A1(g10438A));
NAND2_X1 U_g10479A (.ZN(g10479A),.A2(I16060A),.A1(I16059A));
NAND3_X1 U_g8737A (.ZN(g8737A),.A3(g8688A),.A2(FE_OFN200_g4921A),.A1(g1975A));
NAND2_X1 U_g5942A (.ZN(g5942A),.A2(I9576A),.A1(I9575A));
NAND2_X1 U_g10478A (.ZN(g10478A),.A2(I16053A),.A1(I16052A));
NAND2_X1 U_I12004A (.ZN(I12004A),.A2(I12002A),.A1(g153A));
NAND2_X1 U_I4911A (.ZN(I4911A),.A2(I4910A),.A1(g386A));
NAND2_X1 U_I11914A (.ZN(I11914A),.A2(g1494A),.A1(g5803A));
NAND2_X1 U_g7960A (.ZN(g7960A),.A2(g5573A),.A1(g7409A));
NAND2_X1 U_I5295A (.ZN(I5295A),.A2(g798A),.A1(g794A));
NAND2_X1 U_I12106A (.ZN(I12106A),.A2(g135A),.A1(g6042A));
NAND2_X1 U_I8728A (.ZN(I8728A),.A2(g1117A),.A1(g4605A));
NAND2_X1 U_g3681A (.ZN(g3681A),.A2(I6838A),.A1(I6837A));
NAND2_X1 U_I11907A (.ZN(I11907A),.A2(g1474A),.A1(g5838A));
NAND2_X1 U_I13907A (.ZN(I13907A),.A2(g1432A),.A1(g8265A));
NAND2_X1 U_I8730A (.ZN(I8730A),.A2(I8728A),.A1(g1117A));
NAND2_X1 U_g8551A (.ZN(g8551A),.A2(g8390A),.A1(g3967A));
NAND2_X1 U_I4980A (.ZN(I4980A),.A2(I4978A),.A1(g333A));
NAND2_X1 U_g2961A (.ZN(g2961A),.A2(I6178A),.A1(I6177A));
NAND2_X1 U_g6019A (.ZN(g6019A),.A2(FE_OFN200_g4921A),.A1(g617A));
NAND2_X1 U_I16016A (.ZN(I16016A),.A2(I16015A),.A1(g10441A));
NAND2_X1 U_I11935A (.ZN(I11935A),.A2(g1458A),.A1(g5857A));
NAND2_X1 U_I8678A (.ZN(I8678A),.A2(I8676A),.A1(g1027A));
NAND2_X1 U_I17051A (.ZN(I17051A),.A2(g11249A),.A1(g10923A));
NAND2_X1 U_g4482A (.ZN(g4482A),.A2(I7865A),.A1(I7864A));
NAND2_X1 U_g7592A (.ZN(g7592A),.A2(I12108A),.A1(I12107A));
NAND2_X1 U_g3460A (.ZN(g3460A),.A2(I6666A),.A1(I6665A));
NAND4_X1 U_g7932A (.ZN(g7932A),.A4(FE_OFN96_g2169A),.A3(FE_OFN91_g2172A),.A2(FE_OFN80_g2175A),.A1(g6941A));
NAND2_X1 U_g7624A (.ZN(g7624A),.A2(I12216A),.A1(I12215A));
NAND4_X1 U_g7953A (.ZN(g7953A),.A4(g7550A),.A3(g7562A),.A2(g7574A),.A1(g6941A));
NAND2_X1 U_g8414A (.ZN(g8414A),.A2(I13554A),.A1(I13553A));
NAND2_X1 U_I6168A (.ZN(I6168A),.A2(I6166A),.A1(g153A));
NAND2_X1 U_I5229A (.ZN(I5229A),.A2(g148A),.A1(g182A));
NAND2_X1 U_I6772A (.ZN(I6772A),.A2(I6770A),.A1(g382A));
NAND2_X1 U_I16030A (.ZN(I16030A),.A2(g10430A),.A1(g829A));
NAND2_X1 U_I13284A (.ZN(I13284A),.A2(I13283A),.A1(g1927A));
NAND2_X1 U_I16065A (.ZN(I16065A),.A2(FE_OFN237_g1806A),.A1(g10428A));
NAND2_X1 U_g2947A (.ZN(g2947A),.A2(I6138A),.A1(I6137A));
NAND2_X1 U_I7321A (.ZN(I7321A),.A2(g1231A),.A1(g3047A));
NAND2_X1 U_g2437A (.ZN(g2437A),.A2(I5530A),.A1(I5529A));
NAND2_X1 U_g2102A (.ZN(g2102A),.A2(I4956A),.A1(I4955A));
NAND2_X1 U_I17282A (.ZN(I17282A),.A2(I17281A),.A1(g11221A));
NAND2_X1 U_I5620A (.ZN(I5620A),.A2(I5618A),.A1(FE_OFN247_g1771A));
NAND2_X1 U_I8664A (.ZN(I8664A),.A2(I8662A),.A1(g476A));
NAND2_X1 U_g7524A (.ZN(g7524A),.A2(I11916A),.A1(I11915A));
NAND2_X1 U_g7717A (.ZN(g7717A),.A2(g1950A),.A1(g6863A));
NAND2_X1 U_I16467A (.ZN(I16467A),.A2(g10518A),.A1(g10716A));
NAND2_X1 U_I4972A (.ZN(I4972A),.A2(I4971A),.A1(g991A));
NAND2_X1 U_I13554A (.ZN(I13554A),.A2(I13552A),.A1(g8262A));
NAND2_X1 U_I16037A (.ZN(I16037A),.A2(FE_OFN252_g1791A),.A1(g10363A));
NAND2_X1 U_g8302A (.ZN(g8302A),.A2(I13274A),.A1(I13273A));
NAND2_X1 U_I4943A (.ZN(I4943A),.A2(I4941A),.A1(g324A));
NAND2_X1 U_I5485A (.ZN(I5485A),.A2(I5484A),.A1(g1250A));
NAND2_X1 U_g5527A (.ZN(g5527A),.A2(g4749A),.A1(g3978A));
NAND2_X1 U_I10509A (.ZN(I10509A),.A2(I10507A),.A1(g786A));
NAND2_X1 U_g7599A (.ZN(g7599A),.A2(I12145A),.A1(I12144A));
NAND2_X1 U_I10508A (.ZN(I10508A),.A2(I10507A),.A1(g6221A));
NAND2_X1 U_I6126A (.ZN(I6126A),.A2(I6124A),.A1(g1419A));
NAND2_X1 U_I8671A (.ZN(I8671A),.A2(I8669A),.A1(g814A));
NAND2_X1 U_I6760A (.ZN(I6760A),.A2(g1448A),.A1(g2943A));
NAND2_X1 U_g3626A (.ZN(g3626A),.A2(I6779A),.A1(I6778A));
NAND2_X1 U_I11973A (.ZN(I11973A),.A2(g1462A),.A1(g5852A));
NAND2_X1 U_g2389A (.ZN(g2389A),.A2(I5470A),.A1(I5469A));
NAND2_X1 U_I15617A (.ZN(I15617A),.A2(I15615A),.A1(g10153A));
NAND2_X1 U_g5277A (.ZN(g5277A),.A2(g4538A),.A1(g3734A));
NAND2_X1 U_I5005A (.ZN(I5005A),.A2(g312A),.A1(g421A));
NAND2_X1 U_I6779A (.ZN(I6779A),.A2(I6777A),.A1(g650A));
NAND2_X1 U_I6665A (.ZN(I6665A),.A2(I6664A),.A1(g2792A));
NAND2_X1 U_I8589A (.ZN(I8589A),.A2(g501A),.A1(g4251A));
NAND2_X1 U_g8412A (.ZN(g8412A),.A2(I13546A),.A1(I13545A));
NAND2_X1 U_g2963A (.ZN(g2963A),.A2(I6188A),.A1(I6187A));
NAND2_X1 U_I12045A (.ZN(I12045A),.A2(g1486A),.A1(g5814A));
NAND2_X1 U_I16053A (.ZN(I16053A),.A2(I16051A),.A1(g10434A));
NAND2_X1 U_g2109A (.ZN(g2109A),.A2(I4997A),.A1(I4996A));
NAND2_X1 U_g11418A (.ZN(g11418A),.A2(I17307A),.A1(I17306A));
NAND2_X1 U_I13539A (.ZN(I13539A),.A2(I13537A),.A1(g8157A));
NAND2_X1 U_g10475A (.ZN(g10475A),.A2(I16032A),.A1(I16031A));
NAND2_X1 U_I5324A (.ZN(I5324A),.A2(I5323A),.A1(g1336A));
NAND2_X1 U_I13538A (.ZN(I13538A),.A2(I13537A),.A1(g658A));
NAND2_X1 U_I5469A (.ZN(I5469A),.A2(I5468A),.A1(g1245A));
NAND2_X1 U_I5540A (.ZN(I5540A),.A2(I5538A),.A1(g1023A));
NAND2_X1 U_I17505A (.ZN(I17505A),.A2(I17503A),.A1(g5269A));
NAND2_X1 U_I11241A (.ZN(I11241A),.A2(g790A),.A1(g6760A));
NAND2_X1 U_I8803A (.ZN(I8803A),.A2(g1113A),.A1(g4677A));
NAND2_X1 U_I12061A (.ZN(I12061A),.A2(I12060A),.A1(g5824A));
NAND2_X1 U_I8780A (.ZN(I8780A),.A2(I8778A),.A1(g1137A));
NAND3_X1 U_g8745A (.ZN(g8745A),.A3(I9265A),.A2(g47A),.A1(g8617A));
NAND2_X1 U_I4979A (.ZN(I4979A),.A2(I4978A),.A1(g411A));
NAND2_X1 U_g8109A (.ZN(g8109A),.A2(I11360A),.A1(g48A));
NAND2_X1 U_g8309A (.ZN(g8309A),.A2(I13309A),.A1(I13308A));
NAND2_X1 U_g6758A (.ZN(g6758A),.A2(I10771A),.A1(I10770A));
NAND2_X1 U_I16009A (.ZN(I16009A),.A2(I16007A),.A1(FE_OFN236_g1776A));
NAND2_X1 U_I15616A (.ZN(I15616A),.A2(I15615A),.A1(g10043A));
NAND2_X1 U_I8662A (.ZN(I8662A),.A2(g476A),.A1(g4286A));
NAND2_X1 U_I16008A (.ZN(I16008A),.A2(I16007A),.A1(g10434A));
NAND2_X1 U_I13515A (.ZN(I13515A),.A2(I13513A),.A1(g8248A));
NAND2_X1 U_I13991A (.ZN(I13991A),.A2(I13990A),.A1(g622A));
NAND2_X1 U_g11276A (.ZN(g11276A),.A2(I17053A),.A1(I17052A));
NAND2_X1 U_I15900A (.ZN(I15900A),.A2(I15898A),.A1(g10359A));
NAND2_X1 U_g2419A (.ZN(g2419A),.A2(I5502A),.A1(I5501A));
NAND2_X1 U_I16074A (.ZN(I16074A),.A2(I16072A),.A1(g10438A));
NAND2_X1 U_I10769A (.ZN(I10769A),.A2(FE_OFN251_g1801A),.A1(g5944A));
NAND2_X1 U_I7323A (.ZN(I7323A),.A2(I7321A),.A1(g1231A));
NAND2_X1 U_g7978A (.ZN(g7978A),.A2(g736A),.A1(g7697A));
NAND2_X1 U_I7875A (.ZN(I7875A),.A2(g810A),.A1(g4109A));
NAND2_X1 U_I8562A (.ZN(I8562A),.A2(I8561A),.A1(g4227A));
NAND2_X1 U_I15892A (.ZN(I15892A),.A2(I15890A),.A1(g10285A));
NAND2_X1 U_g3771A (.ZN(g3771A),.A2(I6990A),.A1(I6989A));
NAND2_X1 U_I8605A (.ZN(I8605A),.A2(I8604A),.A1(g4259A));
NAND2_X1 U_g10153A (.ZN(g10153A),.A2(I15453A),.A1(I15452A));
NAND2_X1 U_g5295A (.ZN(g5295A),.A2(I8763A),.A1(I8762A));
NAND2_X1 U_I8751A (.ZN(I8751A),.A2(I8750A),.A1(g4613A));
NAND2_X1 U_I15907A (.ZN(I15907A),.A2(I15906A),.A1(g6899A));
NAND2_X1 U_I5136A (.ZN(I5136A),.A2(I5135A),.A1(g521A));
NAND2_X1 U_I11263A (.ZN(I11263A),.A2(I11261A),.A1(g826A));
NAND2_X1 U_I14204A (.ZN(I14204A),.A2(I14202A),.A1(g591A));
NAND2_X1 U_g8881A (.ZN(g8881A),.A2(I14211A),.A1(I14210A));
NAND2_X1 U_g2105A (.ZN(g2105A),.A2(I4973A),.A1(I4972A));
NAND3_X1 U_g5557A (.ZN(g5557A),.A3(g3011A),.A2(g3071A),.A1(g4538A));
NAND2_X1 U_I5230A (.ZN(I5230A),.A2(I5229A),.A1(g182A));
NAND2_X1 U_I8669A (.ZN(I8669A),.A2(g814A),.A1(g4831A));
NAND2_X1 U_g10474A (.ZN(g10474A),.A2(I16025A),.A1(I16024A));
NAND2_X1 U_I8772A (.ZN(I8772A),.A2(I8770A),.A1(g1133A));
NAND2_X1 U_g2445A (.ZN(g2445A),.A2(I5540A),.A1(I5539A));
NAND2_X1 U_g8006A (.ZN(g8006A),.A2(g7717A),.A1(g5552A));
NAND2_X1 U_I10932A (.ZN(I10932A),.A2(I10930A),.A1(g5555A));
NAND2_X1 U_I17504A (.ZN(I17504A),.A2(I17503A),.A1(g11430A));
NAND2_X1 U_I5137A (.ZN(I5137A),.A2(I5135A),.A1(g525A));
NAND2_X1 U_g8305A (.ZN(g8305A),.A2(I13285A),.A1(I13284A));
NAND2_X1 U_I5891A (.ZN(I5891A),.A2(g2057A),.A1(g750A));
NAND2_X1 U_I13273A (.ZN(I13273A),.A2(I13272A),.A1(g1918A));
NAND2_X1 U_I8480A (.ZN(I8480A),.A2(I8479A),.A1(g4455A));
NAND2_X2 U_g4144A (.ZN(g4144A),.A2(g109A),.A1(g2160A));
NAND2_X1 U_I15906A (.ZN(I15906A),.A2(g10302A),.A1(g6899A));
NAND2_X1 U_I5342A (.ZN(I5342A),.A2(I5341A),.A1(g315A));
NAND2_X1 U_I13514A (.ZN(I13514A),.A2(I13513A),.A1(g686A));
NAND2_X1 U_g8407A (.ZN(g8407A),.A2(I13523A),.A1(I13522A));
NAND2_X1 U_g4088A (.ZN(g4088A),.A2(I7225A),.A1(I7224A));
NAND2_X1 U_g4488A (.ZN(g4488A),.A2(I7877A),.A1(I7876A));
NAND2_X1 U_g7598A (.ZN(g7598A),.A2(I12138A),.A1(I12137A));
NAND3_X1 U_g3222A (.ZN(g3222A),.A3(g1834A),.A2(g1814A),.A1(g2557A));
NAND2_X1 U_I16052A (.ZN(I16052A),.A2(I16051A),.A1(g837A));
NAND2_X1 U_I12127A (.ZN(I12127A),.A2(I12126A),.A1(g6026A));
NAND2_X1 U_g10483A (.ZN(g10483A),.A2(I16088A),.A1(I16087A));
NAND2_X1 U_g8415A (.ZN(g8415A),.A2(I13561A),.A1(I13560A));
NAND2_X1 U_g11415A (.ZN(g11415A),.A2(I17290A),.A1(I17289A));
NAND2_X1 U_g6573A (.ZN(g6573A),.A2(I10509A),.A1(I10508A));
NAND2_X1 U_I5676A (.ZN(I5676A),.A2(I5675A),.A1(g1218A));
NAND2_X1 U_I6778A (.ZN(I6778A),.A2(I6777A),.A1(g2892A));
NAND2_X1 U_g9413A (.ZN(g9413A),.A2(I14614A),.A1(I14613A));
NAND2_X1 U_I8779A (.ZN(I8779A),.A2(I8778A),.A1(g4630A));
NAND2_X1 U_I5592A (.ZN(I5592A),.A2(I5591A),.A1(g1696A));
NAND4_X1 U_g8502A (.ZN(g8502A),.A4(g8366A),.A3(g591A),.A2(g605A),.A1(g2382A));
NAND2_X1 U_I15609A (.ZN(I15609A),.A2(I15607A),.A1(g10144A));
NAND2_X1 U_I15608A (.ZN(I15608A),.A2(I15607A),.A1(g10149A));
NAND3_X1 U_g3071A (.ZN(g3071A),.A3(g2382A),.A2(g2374A),.A1(g605A));
NAND2_X1 U_g10509A (.ZN(g10509A),.A2(g6023A),.A1(g10436A));
NAND2_X1 U_I17461A (.ZN(I17461A),.A2(I17459A),.A1(g11448A));
NAND2_X1 U_I13506A (.ZN(I13506A),.A2(I13504A),.A1(g8247A));
NAND2_X1 U_I5468A (.ZN(I5468A),.A2(g999A),.A1(g1245A));
NAND2_X1 U_g5219A (.ZN(g5219A),.A2(I8652A),.A1(I8651A));
NAND2_X1 U_I5677A (.ZN(I5677A),.A2(I5675A),.A1(g1223A));
NAND3_X1 U_g8826A (.ZN(g8826A),.A3(g8648A),.A2(g8737A),.A1(g8512A));
NAND2_X1 U_I17393A (.ZN(I17393A),.A2(g11414A),.A1(g11415A));
NAND2_X1 U_I5866A (.ZN(I5866A),.A2(I5865A),.A1(g2107A));
NAND2_X1 U_I12126A (.ZN(I12126A),.A2(g170A),.A1(g6026A));
NAND2_X1 U_I4978A (.ZN(I4978A),.A2(g333A),.A1(g411A));
NAND2_X1 U_g7587A (.ZN(g7587A),.A2(I12087A),.A1(I12086A));
NAND2_X1 U_g5286A (.ZN(g5286A),.A2(I8752A),.A1(I8751A));
NAND2_X1 U_g8308A (.ZN(g8308A),.A2(I13302A),.A1(I13301A));
NAND2_X1 U_I7864A (.ZN(I7864A),.A2(I7863A),.A1(g4099A));
NAND2_X1 U_I11981A (.ZN(I11981A),.A2(I11980A),.A1(g5820A));
NAND2_X1 U_I12060A (.ZN(I12060A),.A2(g1478A),.A1(g5824A));
NAND2_X1 U_g5225A (.ZN(g5225A),.A2(I8664A),.A1(I8663A));
NAND2_X1 U_g11538A (.ZN(g11538A),.A2(I17569A),.A1(I17568A));
NAND2_X1 U_I13767A (.ZN(I13767A),.A2(I13765A),.A1(g8417A));
NAND2_X1 U_g10396A (.ZN(g10396A),.A2(I15908A),.A1(I15907A));
NAND2_X1 U_I11262A (.ZN(I11262A),.A2(I11261A),.A1(g6775A));
NAND2_X1 U_I13990A (.ZN(I13990A),.A2(g8688A),.A1(g622A));
NAND2_X1 U_I6224A (.ZN(I6224A),.A2(g1346A),.A1(g2544A));
NAND2_X1 U_I5867A (.ZN(I5867A),.A2(I5865A),.A1(g2105A));
NAND2_X1 U_g2493A (.ZN(g2493A),.A2(g1840A),.A1(g1834A));
NAND2_X1 U_I5893A (.ZN(I5893A),.A2(I5891A),.A1(g2057A));
NAND3_X1 U_g3062A (.ZN(g3062A),.A3(g611A),.A2(g591A),.A1(g2369A));
NAND2_X1 U_I13521A (.ZN(I13521A),.A2(g8249A),.A1(g695A));
NAND2_X1 U_I5186A (.ZN(I5186A),.A2(I5184A),.A1(g1515A));
NAND2_X1 U_I6771A (.ZN(I6771A),.A2(I6770A),.A1(g3257A));
NAND2_X1 U_I5325A (.ZN(I5325A),.A2(I5323A),.A1(g1341A));
NAND2_X1 U_I17459A (.ZN(I17459A),.A2(g11448A),.A1(g11449A));
NAND2_X1 U_I9557A (.ZN(I9557A),.A2(g782A),.A1(g5598A));
NAND2_X1 U_g11414A (.ZN(g11414A),.A2(I17283A),.A1(I17282A));
NAND2_X1 U_I12067A (.ZN(I12067A),.A2(g139A),.A1(g6045A));
NAND2_X1 U_I12094A (.ZN(I12094A),.A2(I12092A),.A1(g1490A));
NAND2_X1 U_I4964A (.ZN(I4964A),.A2(g330A),.A1(g406A));
NAND2_X1 U_I13272A (.ZN(I13272A),.A2(g8158A),.A1(g1918A));
NAND2_X1 U_I9948A (.ZN(I9948A),.A2(I9946A),.A1(g1796A));
NAND2_X1 U_g10302A (.ZN(g10302A),.A2(I15718A),.A1(I15717A));
NAND2_X1 U_I16332A (.ZN(I16332A),.A2(I16330A),.A1(g4997A));
NAND2_X1 U_I5106A (.ZN(I5106A),.A2(I5104A),.A1(g435A));
NAND2_X1 U_g8847A (.ZN(g8847A),.A2(g8683A),.A1(g8551A));
NAND2_X1 U_g2257A (.ZN(g2257A),.A2(I5284A),.A1(I5283A));
NAND2_X1 U_I12019A (.ZN(I12019A),.A2(g166A),.A1(g6049A));
NAND2_X1 U_I15441A (.ZN(I15441A),.A2(g10007A),.A1(g10013A));
NAND2_X1 U_I11997A (.ZN(I11997A),.A2(I11995A),.A1(g127A));
NAND2_X1 U_I8739A (.ZN(I8739A),.A2(I8738A),.A1(g4607A));
NAND2_X1 U_I5461A (.ZN(I5461A),.A2(I5459A),.A1(g1003A));
NAND2_X1 U_I13766A (.ZN(I13766A),.A2(I13765A),.A1(g731A));
NAND2_X1 U_I8479A (.ZN(I8479A),.A2(g3530A),.A1(g4455A));
NAND2_X1 U_I17295A (.ZN(I17295A),.A2(g11227A),.A1(g11229A));
NAND2_X1 U_I14271A (.ZN(I14271A),.A2(I14270A),.A1(g8840A));
NAND2_X1 U_I4971A (.ZN(I4971A),.A2(g995A),.A1(g991A));
NAND2_X1 U_g8301A (.ZN(g8301A),.A2(I13267A),.A1(I13266A));
NAND2_X1 U_I6110A (.ZN(I6110A),.A2(I6109A),.A1(g2205A));
NAND2_X1 U_g10482A (.ZN(g10482A),.A2(I16081A),.A1(I16080A));
NAND2_X1 U_g10779A (.ZN(g10779A),.A2(I16469A),.A1(I16468A));
NAND2_X1 U_I6762A (.ZN(I6762A),.A2(I6760A),.A1(g1448A));
NAND2_X1 U_I17289A (.ZN(I17289A),.A2(I17288A),.A1(g11225A));
NAND2_X1 U_I5315A (.ZN(I5315A),.A2(g1027A),.A1(g1032A));
NAND2_X1 U_I17288A (.ZN(I17288A),.A2(g11223A),.A1(g11225A));
NAND2_X1 U_I13859A (.ZN(I13859A),.A2(I13857A),.A1(g1448A));
NAND2_X1 U_g7548A (.ZN(g7548A),.A2(I11982A),.A1(I11981A));
NAND2_X1 U_I13858A (.ZN(I13858A),.A2(I13857A),.A1(g8270A));
NAND2_X1 U_I11996A (.ZN(I11996A),.A2(I11995A),.A1(g6035A));
NAND3_X1 U_g8743A (.ZN(g8743A),.A3(I9265A),.A2(I9273A),.A1(g8617A));
NAND2_X1 U_I5880A (.ZN(I5880A),.A2(I5878A),.A1(g2115A));
NAND2_X1 U_g10513A (.ZN(g10513A),.A2(g5345A),.A1(g10441A));
NAND2_X1 U_g8411A (.ZN(g8411A),.A2(I13539A),.A1(I13538A));
NAND2_X1 U_I8626A (.ZN(I8626A),.A2(I8624A),.A1(g511A));
NAND2_X1 U_g10505A (.ZN(g10505A),.A2(g5938A),.A1(g10432A));
NAND2_X1 U_I5612A (.ZN(I5612A),.A2(I5611A),.A1(g1280A));
NAND2_X1 U_g4821A (.ZN(g4821A),.A2(I8180A),.A1(I8179A));
NAND2_X1 U_I12076A (.ZN(I12076A),.A2(I12074A),.A1(g174A));
NAND2_X1 U_I12085A (.ZN(I12085A),.A2(g1470A),.A1(g5842A));
NAND2_X1 U_g7567A (.ZN(g7567A),.A2(I12021A),.A1(I12020A));
NAND2_X1 U_I5128A (.ZN(I5128A),.A2(I5126A),.A1(g1389A));
NAND2_X1 U_I6489A (.ZN(I6489A),.A2(I6487A),.A1(g1227A));
NAND2_X1 U_g7593A (.ZN(g7593A),.A2(I12115A),.A1(I12114A));
NAND2_X1 U_I8778A (.ZN(I8778A),.A2(g1137A),.A1(g4630A));
NAND2_X1 U_g10149A (.ZN(g10149A),.A2(I15443A),.A1(I15442A));
NAND2_X1 U_I13902A (.ZN(I13902A),.A2(I13900A),.A1(g1428A));
NAND2_X1 U_I13301A (.ZN(I13301A),.A2(I13300A),.A1(g1936A));
NAND2_X1 U_g3215A (.ZN(g3215A),.A2(g1822A),.A1(g2564A));
NAND4_X1 U_g7996A (.ZN(g7996A),.A4(FE_OFN96_g2169A),.A3(g7562A),.A2(g7574A),.A1(FE_OFN88_g2178A));
NAND2_X1 U_I4985A (.ZN(I4985A),.A2(g1003A),.A1(g999A));
NAND2_X1 U_I14444A (.ZN(I14444A),.A2(I14442A),.A1(g1834A));
NAND4_X1 U_g8000A (.ZN(g8000A),.A4(g7550A),.A3(g7562A),.A2(g7574A),.A1(FE_OFN88_g2178A));
NAND2_X1 U_I5166A (.ZN(I5166A),.A2(I5164A),.A1(g1499A));
NAND2_X1 U_I17460A (.ZN(I17460A),.A2(I17459A),.A1(g11449A));
NAND2_X1 U_g3008A (.ZN(g3008A),.A2(g878A),.A1(g2444A));
NAND2_X1 U_I6836A (.ZN(I6836A),.A2(g806A),.A1(g3287A));
NAND2_X1 U_I5529A (.ZN(I5529A),.A2(I5528A),.A1(g1265A));
NAND2_X1 U_g10229A (.ZN(g10229A),.A2(I15609A),.A1(I15608A));
NAND2_X1 U_I13661A (.ZN(I13661A),.A2(I13659A),.A1(g8322A));
NAND2_X1 U_I13895A (.ZN(I13895A),.A2(I13893A),.A1(g1436A));
NAND2_X1 U_g2303A (.ZN(g2303A),.A2(I5343A),.A1(I5342A));
NAND2_X1 U_I12039A (.ZN(I12039A),.A2(I12038A),.A1(g5847A));
NAND2_X1 U_g5592A (.ZN(g5592A),.A2(I9008A),.A1(I9007A));
NAND2_X1 U_I12038A (.ZN(I12038A),.A2(g1466A),.A1(g5847A));
NAND2_X1 U_g3322A (.ZN(g3322A),.A2(I6489A),.A1(I6488A));
NAND2_X1 U_I8561A (.ZN(I8561A),.A2(g491A),.A1(g4227A));
NAND2_X1 U_I8527A (.ZN(I8527A),.A2(g481A),.A1(g4879A));
NAND2_X1 U_I12143A (.ZN(I12143A),.A2(g158A),.A1(g6000A));
NAND2_X1 U_I5619A (.ZN(I5619A),.A2(I5618A),.A1(g1766A));
NAND2_X1 U_g10386A (.ZN(g10386A),.A2(I15880A),.A1(I15879A));
NAND2_X1 U_I11980A (.ZN(I11980A),.A2(g1482A),.A1(g5820A));
NAND2_X1 U_I6837A (.ZN(I6837A),.A2(I6836A),.A1(g3287A));
NAND2_X1 U_I4973A (.ZN(I4973A),.A2(I4971A),.A1(g995A));
NAND2_X1 U_I13888A (.ZN(I13888A),.A2(I13886A),.A1(g1440A));
NAND2_X1 U_g7558A (.ZN(g7558A),.A2(I12004A),.A1(I12003A));
NAND2_X1 U_I17494A (.ZN(I17494A),.A2(I17492A),.A1(g3623A));
NAND2_X1 U_g11491A (.ZN(g11491A),.A2(I17494A),.A1(I17493A));
NAND2_X1 U_I16045A (.ZN(I16045A),.A2(I16044A),.A1(g833A));
NAND2_X1 U_I7684A (.ZN(I7684A),.A2(I7683A),.A1(g1023A));
NAND2_X1 U_g4130A (.ZN(g4130A),.A2(g2518A),.A1(FE_OFN352_g109A));
NAND2_X1 U_I8771A (.ZN(I8771A),.A2(I8770A),.A1(g4619A));
NAND2_X1 U_I13546A (.ZN(I13546A),.A2(I13544A),.A1(g8259A));
NAND2_X1 U_I13089A (.ZN(I13089A),.A2(g1840A),.A1(g8006A));
NAND2_X1 U_g2117A (.ZN(g2117A),.A2(I5025A),.A1(I5024A));
NAND2_X1 U_g5119A (.ZN(g5119A),.A2(I8515A),.A1(I8514A));
NAND2_X1 U_g5319A (.ZN(g5319A),.A2(I8805A),.A1(I8804A));
NAND2_X1 U_I15899A (.ZN(I15899A),.A2(I15898A),.A1(g857A));
NAND2_X1 U_I5606A (.ZN(I5606A),.A2(I5604A),.A1(g1153A));
NAND2_X1 U_I15898A (.ZN(I15898A),.A2(g10359A),.A1(g857A));
NAND2_X1 U_I16032A (.ZN(I16032A),.A2(I16030A),.A1(g10430A));
NAND2_X1 U_I17401A (.ZN(I17401A),.A2(I17400A),.A1(g11418A));
NAND2_X1 U_I13659A (.ZN(I13659A),.A2(g8322A),.A1(g1945A));
NAND2_X1 U_I8738A (.ZN(I8738A),.A2(g1121A),.A1(g4607A));
NAND2_X1 U_I13250A (.ZN(I13250A),.A2(I13248A),.A1(g8148A));
NAND2_X1 U_I15718A (.ZN(I15718A),.A2(I15716A),.A1(g10229A));
NAND2_X1 U_I9008A (.ZN(I9008A),.A2(I9006A),.A1(FE_OFN252_g1791A));
NAND2_X1 U_I6176A (.ZN(I6176A),.A2(g197A),.A1(g2177A));
NAND2_X1 U_I7865A (.ZN(I7865A),.A2(I7863A),.A1(g774A));
NAND2_X1 U_g5274A (.ZN(g5274A),.A2(I8730A),.A1(I8729A));
NAND2_X1 U_I5341A (.ZN(I5341A),.A2(g426A),.A1(g315A));
NAND2_X1 U_I17305A (.ZN(I17305A),.A2(g11231A),.A1(g11232A));
NAND2_X1 U_I17053A (.ZN(I17053A),.A2(I17051A),.A1(g11249A));
NAND2_X1 U_g5125A (.ZN(g5125A),.A2(I8529A),.A1(I8528A));
NAND2_X1 U_I12216A (.ZN(I12216A),.A2(I12214A),.A1(g2518A));
NAND2_X1 U_I6225A (.ZN(I6225A),.A2(I6224A),.A1(g2544A));
NAND2_X1 U_I5879A (.ZN(I5879A),.A2(I5878A),.A1(g2120A));
NAND2_X1 U_g3221A (.ZN(g3221A),.A2(g2564A),.A1(g1834A));
NAND2_X1 U_I14270A (.ZN(I14270A),.A2(g1822A),.A1(g8840A));
NAND2_X1 U_I6124A (.ZN(I6124A),.A2(g1419A),.A1(g2215A));
NAND2_X1 U_I6324A (.ZN(I6324A),.A2(I6322A),.A1(g1864A));
NAND2_X1 U_I13867A (.ZN(I13867A),.A2(g1403A),.A1(g8264A));
NAND2_X1 U_I13894A (.ZN(I13894A),.A2(I13893A),.A1(g8266A));
NAND2_X1 U_I6469A (.ZN(I6469A),.A2(I6467A),.A1(g2479A));
NAND2_X1 U_I8663A (.ZN(I8663A),.A2(I8662A),.A1(g4286A));
NAND2_X1 U_g7523A (.ZN(g7523A),.A2(I11909A),.A1(I11908A));
NAND2_X1 U_I6177A (.ZN(I6177A),.A2(I6176A),.A1(g2177A));
NAND2_X1 U_g5187A (.ZN(g5187A),.A2(I8591A),.A1(I8590A));
NAND2_X1 U_I6287A (.ZN(I6287A),.A2(g981A),.A1(g2091A));
NAND2_X1 U_I8762A (.ZN(I8762A),.A2(I8761A),.A1(g4616A));
NAND2_X1 U_I15871A (.ZN(I15871A),.A2(I15870A),.A1(g10291A));
NAND3_X1 U_g8840A (.ZN(g8840A),.A3(g8551A),.A2(g8541A),.A1(g8542A));
NAND2_X1 U_g2250A (.ZN(g2250A),.A2(I5265A),.A1(I5264A));
NAND2_X1 U_I8590A (.ZN(I8590A),.A2(I8589A),.A1(g4251A));
NAND2_X1 U_I6199A (.ZN(I6199A),.A2(g766A),.A1(g2525A));
NAND2_X1 U_I14218A (.ZN(I14218A),.A2(I14216A),.A1(g605A));
NAND2_X1 U_g8190A (.ZN(g8190A),.A2(g7978A),.A1(g6027A));
NAND2_X1 U_I5284A (.ZN(I5284A),.A2(I5282A),.A1(g762A));
NAND2_X1 U_I17485A (.ZN(I17485A),.A2(g11474A),.A1(g11233A));
NAND2_X1 U_I4965A (.ZN(I4965A),.A2(I4964A),.A1(g406A));
NAND2_X1 U_I5591A (.ZN(I5591A),.A2(g1703A),.A1(g1696A));
NAND2_X1 U_g8501A (.ZN(g8501A),.A2(g8366A),.A1(g3760A));
NAND2_X1 U_I15451A (.ZN(I15451A),.A2(g10019A),.A1(g10025A));
NAND2_X1 U_g8942A (.ZN(g8942A),.A2(FE_OFN200_g4921A),.A1(g8823A));
NAND2_X1 U_I13877A (.ZN(I13877A),.A2(I13876A),.A1(g8269A));
NAND2_X1 U_g7269A (.ZN(g7269A),.A2(I11510A),.A1(I11509A));
NAND2_X1 U_I4996A (.ZN(I4996A),.A2(I4995A),.A1(g416A));
NAND2_X1 U_I6144A (.ZN(I6144A),.A2(I6143A),.A1(g1976A));
NAND2_X1 U_I17567A (.ZN(I17567A),.A2(g1610A),.A1(g11496A));
NAND2_X1 U_g7572A (.ZN(g7572A),.A2(I12040A),.A1(I12039A));
NAND2_X1 U_I6207A (.ZN(I6207A),.A2(g802A),.A1(g5188A));
NAND2_X1 U_I14277A (.ZN(I14277A),.A2(g1828A),.A1(g8847A));
NAND2_X1 U_I16059A (.ZN(I16059A),.A2(I16058A),.A1(g841A));
NAND2_X1 U_I16025A (.ZN(I16025A),.A2(I16023A),.A1(FE_OFN253_g1786A));
NAND2_X1 U_I8563A (.ZN(I8563A),.A2(I8561A),.A1(g491A));
NAND2_X1 U_g3524A (.ZN(g3524A),.A2(g3221A),.A1(g3209A));
NAND2_X1 U_I16058A (.ZN(I16058A),.A2(g10441A),.A1(g841A));
NAND2_X1 U_I5204A (.ZN(I5204A),.A2(I5202A),.A1(g374A));
NAND2_X1 U_I6488A (.ZN(I6488A),.A2(I6487A),.A1(g2306A));
NAND4_X1 U_g3818A (.ZN(g3818A),.A4(g3003A),.A3(g2310A),.A2(g3071A),.A1(g3056A));
NAND2_X1 U_I16044A (.ZN(I16044A),.A2(g10432A),.A1(g833A));
NAND2_X1 U_g3717A (.ZN(g3717A),.A2(I6881A),.A1(I6880A));
NAND2_X1 U_I13077A (.ZN(I13077A),.A2(I13076A),.A1(g1872A));
NAND2_X1 U_g10043A (.ZN(g10043A),.A2(I15258A),.A1(I15257A));
NAND2_X1 U_I11280A (.ZN(I11280A),.A2(I11278A),.A1(g6485A));
NAND2_X1 U_I6825A (.ZN(I6825A),.A2(g770A),.A1(g3281A));
NAND2_X1 U_I4997A (.ZN(I4997A),.A2(I4995A),.A1(g309A));
NAND2_X1 U_I13300A (.ZN(I13300A),.A2(g8162A),.A1(g1936A));
NAND2_X1 U_I5323A (.ZN(I5323A),.A2(g1341A),.A1(g1336A));
NAND2_X1 U_I6136A (.ZN(I6136A),.A2(g378A),.A1(g2496A));
NAND2_X1 U_g5935A (.ZN(g5935A),.A2(I9559A),.A1(I9558A));
NAND2_X1 U_I5528A (.ZN(I5528A),.A2(g1015A),.A1(g1265A));
NAND2_X1 U_I6806A (.ZN(I6806A),.A2(I6805A),.A1(g3268A));
NAND2_X1 U_I5530A (.ZN(I5530A),.A2(I5528A),.A1(g1015A));
NAND2_X1 U_g10886A (.ZN(g10886A),.A2(g10805A),.A1(g10807A));
NAND2_X1 U_g3106A (.ZN(g3106A),.A2(I6324A),.A1(I6323A));
NAND2_X1 U_I13876A (.ZN(I13876A),.A2(g1444A),.A1(g8269A));
NAND2_X1 U_I6322A (.ZN(I6322A),.A2(g1864A),.A1(g2050A));
NAND2_X1 U_g3061A (.ZN(g3061A),.A2(g2374A),.A1(g611A));
NAND2_X1 U_g2439A (.ZN(g2439A),.A2(g1828A),.A1(g1814A));
NAND4_X1 U_g7947A (.ZN(g7947A),.A4(g7550A),.A3(FE_OFN91_g2172A),.A2(g7574A),.A1(g6941A));
NAND2_X1 U_I9576A (.ZN(I9576A),.A2(I9574A),.A1(g818A));
NAND2_X1 U_I13660A (.ZN(I13660A),.A2(I13659A),.A1(g1945A));
NAND2_X1 U_g3200A (.ZN(g3200A),.A2(g2061A),.A1(g1822A));
NAND2_X1 U_g4374A (.ZN(g4374A),.A2(I7685A),.A1(I7684A));
NAND2_X1 U_I11916A (.ZN(I11916A),.A2(I11914A),.A1(g1494A));
NAND2_X1 U_I5372A (.ZN(I5372A),.A2(I5371A),.A1(g971A));
NAND2_X1 U_g3003A (.ZN(g3003A),.A2(g2399A),.A1(g599A));
NAND2_X1 U_g8627A (.ZN(g8627A),.A2(I13888A),.A1(I13887A));
NAND2_X1 U_I5618A (.ZN(I5618A),.A2(FE_OFN247_g1771A),.A1(g1766A));
NAND2_X1 U_I6137A (.ZN(I6137A),.A2(I6136A),.A1(g2496A));
NAND2_X1 U_I5343A (.ZN(I5343A),.A2(I5341A),.A1(g426A));
NAND2_X1 U_I5282A (.ZN(I5282A),.A2(g762A),.A1(g758A));
NAND2_X1 U_I13307A (.ZN(I13307A),.A2(g617A),.A1(g8190A));
NAND2_X1 U_I13076A (.ZN(I13076A),.A2(g7963A),.A1(g1872A));
NAND2_X1 U_I6807A (.ZN(I6807A),.A2(I6805A),.A1(g471A));
NAND2_X1 U_I11243A (.ZN(I11243A),.A2(I11241A),.A1(g790A));
NAND2_X1 U_I17585A (.ZN(I17585A),.A2(I17584A),.A1(g11217A));
NAND2_X1 U_I12137A (.ZN(I12137A),.A2(I12136A),.A1(g6038A));
NAND2_X1 U_I7564A (.ZN(I7564A),.A2(I7562A),.A1(g654A));
NAND2_X1 U_g2970A (.ZN(g2970A),.A2(I6201A),.A1(I6200A));
NAND2_X1 U_g10144A (.ZN(g10144A),.A2(I15432A),.A1(I15431A));
NAND2_X1 U_I8788A (.ZN(I8788A),.A2(I8786A),.A1(g1141A));
NAND2_X1 U_g7054A (.ZN(g7054A),.A2(I11243A),.A1(I11242A));
NAND2_X1 U_I17052A (.ZN(I17052A),.A2(I17051A),.A1(g10923A));
NAND2_X1 U_g2120A (.ZN(g2120A),.A2(I5036A),.A1(I5035A));
NAND2_X1 U_g8616A (.ZN(g8616A),.A2(I13869A),.A1(I13868A));
NAND2_X1 U_I5202A (.ZN(I5202A),.A2(g374A),.A1(g369A));
NAND2_X1 U_I16088A (.ZN(I16088A),.A2(I16086A),.A1(g10430A));
NAND2_X1 U_I16024A (.ZN(I16024A),.A2(I16023A),.A1(g10438A));
NAND2_X1 U_g11490A (.ZN(g11490A),.A2(I17487A),.A1(I17486A));
NAND2_X1 U_I5518A (.ZN(I5518A),.A2(I5516A),.A1(g1019A));
NAND3_X1 U_g5118A (.ZN(g5118A),.A3(g4073A),.A2(g4806A),.A1(g2439A));
NAND2_X1 U_I12021A (.ZN(I12021A),.A2(I12019A),.A1(g166A));
NOR2_X1 U_g6392A (.ZN(g6392A),.A2(g5938A),.A1(g5859A));
NOR2_X1 U_g5938A (.ZN(g5938A),.A2(FE_OFN349_I6424A),.A1(g2273A));
NOR2_X1 U_g2478A (.ZN(g2478A),.A2(g1737A),.A1(g1610A));
NOR4_X1 U_g4278A (.ZN(g4278A),.A4(g3776A),.A3(FE_OFN254_g461A),.A2(FE_OFN248_g466A),.A1(g3800A));
NOR2_X1 U_g10383A (.ZN(g10383A),.A2(g3348A),.A1(I15514A));
NOR2_X1 U_g3118A (.ZN(g3118A),.A2(g2514A),.A1(g2521A));
NOR2_X1 U_g9815A (.ZN(g9815A),.A2(FE_OFN67_g9367A),.A1(FE_OFN68_g9392A));
NOR2_X1 U_g11077A (.ZN(g11077A),.A2(g10971A),.A1(g10970A));
NOR3_X1 U_g3879A (.ZN(g3879A),.A3(g2353A),.A2(g2354A),.A1(g3141A));
NOR2_X1 U_g10285A (.ZN(g10285A),.A2(FE_OFN350_g3121A),.A1(I15287A));
NOR2_X1 U_g11480A (.ZN(g11480A),.A2(g4567A),.A1(g11456A));
NOR2_X1 U_g4076A (.ZN(g4076A),.A2(I5254A),.A1(g1707A));
NOR2_X1 U_g10570A (.ZN(g10570A),.A2(g10324A),.A1(g10485A));
NOR2_X1 U_g10239A (.ZN(g10239A),.A2(I15287A),.A1(g9317A));
NOR2_X1 U_g10594A (.ZN(g10594A),.A2(g10521A),.A1(g10480A));
NOR2_X1 U_g9426A (.ZN(g9426A),.A2(FE_OFN50_g9030A),.A1(FE_OFN54_g9052A));
NOR2_X1 U_g10382A (.ZN(g10382A),.A2(g3348A),.A1(I15507A));
NOR4_X1 U_g4672A (.ZN(g4672A),.A4(g3479A),.A3(g1104A),.A2(g1107A),.A1(g3501A));
NOR2_X1 U_g5360A (.ZN(g5360A),.A2(FE_OFN308_I6424A),.A1(g105A));
NOR4_X1 U_g9387A (.ZN(g9387A),.A4(I14779A),.A3(g9223A),.A2(g9240A),.A1(g9010A));
NOR2_X1 U_g10438A (.ZN(g10438A),.A2(FE_OFN160_I6424A),.A1(I15500A));
NOR4_X1 U_g4613A (.ZN(g4613A),.A4(g1101A),.A3(g1104A),.A2(g3491A),.A1(FE_OFN240_g1110A));
NOR4_X1 U_g9391A (.ZN(g9391A),.A4(I14602A),.A3(FE_OFN39_g9223A),.A2(FE_OFN40_g9240A),.A1(g9010A));
NOR3_X1 U_g4572A (.ZN(g4572A),.A3(g3628A),.A2(g3408A),.A1(g3419A));
NOR3_X1 U_g9757A (.ZN(g9757A),.A3(FE_OFN72_g9292A),.A2(FE_OFN62_g9274A),.A1(FE_OFN32_g9454A));
NOR4_X1 U_g9874A (.ZN(g9874A),.A4(I15033A),.A3(g9579A),.A2(FE_OFN64_g9536A),.A1(g9519A));
NOR2_X1 U_g9654A (.ZN(g9654A),.A2(FE_OFN53_g9173A),.A1(FE_OFN46_g9125A));
NOR4_X1 U_g9880A (.ZN(g9880A),.A4(I15051A),.A3(g9579A),.A2(FE_OFN64_g9536A),.A1(g9751A));
NOR4_X1 U_g4873A (.ZN(g4873A),.A4(g3776A),.A3(FE_OFN254_g461A),.A2(FE_OFN248_g466A),.A1(FE_OFN250_g471A));
NOR2_X1 U_g2807A (.ZN(g2807A),.A2(g3629A),.A1(FE_OFN266_g18A));
NOR2_X1 U_g10441A (.ZN(g10441A),.A2(FE_OFN160_I6424A),.A1(I15510A));
NOR4_X1 U_g4639A (.ZN(g4639A),.A4(g1101A),.A3(g1104A),.A2(g1107A),.A1(g3501A));
NOR2_X1 U_g10435A (.ZN(g10435A),.A2(g3744A),.A1(I15510A));
NOR2_X1 U_g10849A (.ZN(g10849A),.A2(g2459A),.A1(g10739A));
NOR4_X1 U_g9606A (.ZN(g9606A),.A4(FE_OFN48_g9151A),.A3(FE_OFN52_g9173A),.A2(FE_OFN51_g9111A),.A1(FE_OFN45_g9125A));
NOR4_X1 U_g9879A (.ZN(g9879A),.A4(I15048A),.A3(g9563A),.A2(FE_OFN64_g9536A),.A1(g9747A));
NOR2_X1 U_g9506A (.ZN(g9506A),.A2(FE_OFN49_g9030A),.A1(FE_OFN56_g9052A));
NOR2_X1 U_g6155A (.ZN(g6155A),.A2(I5254A),.A1(g4974A));
NOR2_X1 U_g6355A (.ZN(g6355A),.A2(g6023A),.A1(g6032A));
NOR2_X1 U_g9591A (.ZN(g9591A),.A2(FE_OFN47_g9151A),.A1(FE_OFN44_g9125A));
NOR2_X1 U_g10359A (.ZN(g10359A),.A2(FE_OFN308_I6424A),.A1(I15290A));
NOR2_X1 U_g10434A (.ZN(g10434A),.A2(FE_OFN349_I6424A),.A1(I15514A));
NOR2_X1 U_g10291A (.ZN(g10291A),.A2(FE_OFN308_I6424A),.A1(I15287A));
NOR4_X1 U_g4227A (.ZN(g4227A),.A4(g2579A),.A3(FE_OFN254_g461A),.A2(g3793A),.A1(FE_OFN250_g471A));
NOR4_X1 U_g9667A (.ZN(g9667A),.A4(FE_OFN47_g9151A),.A3(FE_OFN52_g9173A),.A2(FE_OFN51_g9111A),.A1(FE_OFN45_g9125A));
NOR2_X1 U_g10563A (.ZN(g10563A),.A2(g10322A),.A1(g10484A));
NOR2_X1 U_g10324A (.ZN(g10324A),.A2(I15365A),.A1(g9317A));
NOR3_X1 U_g4455A (.ZN(g4455A),.A3(g3408A),.A2(g3419A),.A1(g3543A));
NOR4_X1 U_g9878A (.ZN(g9878A),.A4(I15045A),.A3(g9579A),.A2(FE_OFN64_g9536A),.A1(g9754A));
NOR2_X1 U_g10360A (.ZN(g10360A),.A2(FE_OFN350_g3121A),.A1(I15290A));
NOR4_X1 U_g9882A (.ZN(g9882A),.A4(I15057A),.A3(g9563A),.A2(FE_OFN64_g9536A),.A1(g9747A));
NOR4_X1 U_g4605A (.ZN(g4605A),.A4(g1101A),.A3(g3485A),.A2(g1107A),.A1(FE_OFN240_g1110A));
NOR2_X1 U_g10562A (.ZN(g10562A),.A2(g10529A),.A1(g10483A));
NOR2_X1 U_g5780A (.ZN(g5780A),.A2(FE_OFN200_g4921A),.A1(g3092A));
NOR2_X1 U_g10385A (.ZN(g10385A),.A2(g3348A),.A1(I15510A));
NOR4_X1 U_g4601A (.ZN(g4601A),.A4(g3479A),.A3(g1104A),.A2(g1107A),.A1(FE_OFN240_g1110A));
NOR2_X1 U_g5573A (.ZN(g5573A),.A2(g4432A),.A1(g4117A));
NOR2_X1 U_g5999A (.ZN(g5999A),.A2(FE_OFN349_I6424A),.A1(g2271A));
NOR3_X1 U_g9759A (.ZN(g9759A),.A3(FE_OFN71_g9292A),.A2(g9274A),.A1(g9454A));
NOR2_X1 U_g6037A (.ZN(g6037A),.A2(FE_OFN350_g3121A),.A1(g2297A));
NOR2_X1 U_g5034A (.ZN(g5034A),.A2(g3967A),.A1(g3524A));
NOR4_X1 U_g9881A (.ZN(g9881A),.A4(I15054A),.A3(g9579A),.A2(FE_OFN64_g9536A),.A1(g9516A));
NOR3_X1 U_g4276A (.ZN(g4276A),.A3(g2500A),.A2(g3261A),.A1(g4065A));
NOR4_X1 U_g4616A (.ZN(g4616A),.A4(g3479A),.A3(g1104A),.A2(g3491A),.A1(FE_OFN240_g1110A));
NOR2_X1 U_g10363A (.ZN(g10363A),.A2(FE_OFN308_I6424A),.A1(I15365A));
NOR2_X1 U_g2862A (.ZN(g2862A),.A2(g2305A),.A1(g2315A));
NOR3_X1 U_g9758A (.ZN(g9758A),.A3(FE_OFN71_g9292A),.A2(FE_OFN62_g9274A),.A1(FE_OFN32_g9454A));
NOR3_X1 U_g9589A (.ZN(g9589A),.A3(FE_OFN48_g9151A),.A2(FE_OFN52_g9173A),.A1(FE_OFN45_g9125A));
NOR2_X1 U_g9803A (.ZN(g9803A),.A2(g9367A),.A1(FE_OFN69_g9392A));
NOR2_X1 U_g10430A (.ZN(g10430A),.A2(FE_OFN349_I6424A),.A1(I15503A));
NOR2_X1 U_g10362A (.ZN(g10362A),.A2(g3744A),.A1(I15290A));
NOR2_X1 U_g2791A (.ZN(g2791A),.A2(g750A),.A1(g2187A));
NOR4_X1 U_g9605A (.ZN(g9605A),.A4(FE_OFN48_g9151A),.A3(FE_OFN52_g9173A),.A2(FE_OFN51_g9111A),.A1(FE_OFN46_g9125A));
NOR2_X1 U_g10436A (.ZN(g10436A),.A2(FE_OFN349_I6424A),.A1(I15510A));
NOR4_X1 U_g5556A (.ZN(g5556A),.A4(g2031A),.A3(g2299A),.A2(FE_OFN238_g1781A),.A1(g4787A));
NOR4_X1 U_g4286A (.ZN(g4286A),.A4(g2579A),.A3(g3784A),.A2(FE_OFN248_g466A),.A1(g3800A));
NOR2_X1 U_g4974A (.ZN(g4974A),.A2(g3714A),.A1(g4502A));
NOR2_X1 U_g9423A (.ZN(g9423A),.A2(FE_OFN49_g9030A),.A1(FE_OFN54_g9052A));
NOR2_X1 U_g5350A (.ZN(g5350A),.A2(FE_OFN160_I6424A),.A1(g3070A));
NOR4_X1 U_g2459A (.ZN(g2459A),.A4(g1648A),.A3(g1651A),.A2(g1642A),.A1(g1645A));
NOR2_X1 U_g10381A (.ZN(g10381A),.A2(g3348A),.A1(I15503A));
NOR4_X1 U_g4259A (.ZN(g4259A),.A4(g3776A),.A3(g3784A),.A2(g3793A),.A1(FE_OFN250_g471A));
NOR2_X1 U_g10522A (.ZN(g10522A),.A2(g10239A),.A1(g10401A));
NOR2_X1 U_g5392A (.ZN(g5392A),.A2(FE_OFN160_I6424A),.A1(g3086A));
NOR3_X1 U_g4122A (.ZN(g4122A),.A3(g2538A),.A2(g2410A),.A1(g3291A));
NOR2_X1 U_g6023A (.ZN(g6023A),.A2(FE_OFN160_I6424A),.A1(g2275A));
NOR2_X1 U_g3462A (.ZN(g3462A),.A2(g2795A),.A1(g2187A));
NOR4_X1 U_g4218A (.ZN(g4218A),.A4(g3776A),.A3(g3784A),.A2(FE_OFN248_g466A),.A1(FE_OFN250_g471A));
NOR4_X1 U_g4267A (.ZN(g4267A),.A4(g2579A),.A3(FE_OFN254_g461A),.A2(FE_OFN248_g466A),.A1(g3800A));
NOR4_X1 U_g4677A (.ZN(g4677A),.A4(g1101A),.A3(g3485A),.A2(g1107A),.A1(g3501A));
NOR2_X1 U_g9646A (.ZN(g9646A),.A2(FE_OFN47_g9151A),.A1(FE_OFN45_g9125A));
NOR2_X1 U_g2863A (.ZN(g2863A),.A2(g2309A),.A1(g2316A));
NOR2_X1 U_g6032A (.ZN(g6032A),.A2(FE_OFN349_I6424A),.A1(g3008A));
NOR4_X1 U_g9647A (.ZN(g9647A),.A4(FE_OFN48_g9151A),.A3(FE_OFN53_g9173A),.A2(FE_OFN51_g9111A),.A1(FE_OFN46_g9125A));
NOR2_X1 U_g5859A (.ZN(g5859A),.A2(FE_OFN349_I6424A),.A1(g2987A));
NOR2_X1 U_g10433A (.ZN(g10433A),.A2(g3744A),.A1(I15514A));
NOR4_X1 U_g4251A (.ZN(g4251A),.A4(g2579A),.A3(g3784A),.A2(g3793A),.A1(FE_OFN250_g471A));
NOR4_X1 U_g9876A (.ZN(g9876A),.A4(I15054A),.A3(FE_OFN56_g9052A),.A2(FE_OFN280_g9536A),.A1(g9522A));
NOR2_X1 U_g8303A (.ZN(g8303A),.A2(g4811A),.A1(g8209A));
NOR2_X1 U_g10429A (.ZN(g10429A),.A2(g3744A),.A1(I15503A));
NOR2_X1 U_g10428A (.ZN(g10428A),.A2(g3121A),.A1(I15503A));
NOR4_X1 U_g4234A (.ZN(g4234A),.A4(g3776A),.A3(FE_OFN254_g461A),.A2(g3793A),.A1(FE_OFN250_g471A));
NOR4_X1 U_g9877A (.ZN(g9877A),.A4(I15048A),.A3(g9569A),.A2(FE_OFN64_g9536A),.A1(g9512A));
NOR2_X1 U_g5186A (.ZN(g5186A),.A2(FE_OFN223_g4401A),.A1(g2047A));
NOR4_X1 U_g4619A (.ZN(g4619A),.A4(g1101A),.A3(g3485A),.A2(g3491A),.A1(FE_OFN240_g1110A));
NOR2_X1 U_g10432A (.ZN(g10432A),.A2(FE_OFN349_I6424A),.A1(I15507A));
NOR2_X1 U_g5345A (.ZN(g5345A),.A2(FE_OFN350_g3121A),.A1(g2067A));
NOR2_X1 U_g5763A (.ZN(g5763A),.A2(g5345A),.A1(g5350A));
NOR4_X1 U_g4879A (.ZN(g4879A),.A4(g2579A),.A3(g3784A),.A2(FE_OFN248_g466A),.A1(FE_OFN250_g471A));
NOR4_X1 U_g4607A (.ZN(g4607A),.A4(g3479A),.A3(g3485A),.A2(g1107A),.A1(FE_OFN240_g1110A));
NOR2_X1 U_g3107A (.ZN(g3107A),.A2(g2499A),.A1(g2501A));
NOR2_X1 U_g10322A (.ZN(g10322A),.A2(I15500A),.A1(g9317A));
NOR4_X1 U_g4630A (.ZN(g4630A),.A4(g3479A),.A3(g3485A),.A2(g3491A),.A1(FE_OFN240_g1110A));
NOR2_X1 U_g10364A (.ZN(g10364A),.A2(g3744A),.A1(I15507A));
SDFF_X1 U_g1289A (.Q(g1289A),.SE(test_seA),.SI(test_siA),.D(g4556A),.CK(CKA));
SDFF_X1 U_g1882A (.Q(g1882A),.SE(test_seA),.SI(g1289A),.D(g8943A),.CK(CKA));
SDFF_X1 U_g312A (.Q(g312A),.SE(test_seA),.SI(g1882A),.D(g255A),.CK(CKA));
SDFF_X1 U_g452A (.Q(g452A),.SE(test_seA),.SI(g312A),.D(g11257A),.CK(CKA));
SDFF_X1 U_g123A (.Q(g123A),.SE(test_seA),.SI(g452A),.D(g7032A),.CK(CKA));
SDFF_X1 U_g207A (.Q(g207A),.SE(test_seA),.SI(g123A),.D(g6830A),.CK(CKA));
SDFF_X1 U_g713A (.Q(g713A),.SE(test_seA),.SI(g207A),.D(g8920A),.CK(CKA));
SDFF_X1 U_g1153A (.Q(g1153A),.SE(test_seA),.SI(g713A),.D(g4340A),.CK(CKA));
SDFF_X1 U_g1209A (.Q(g1209A),.SE(test_seA),.SI(g1153A),.D(g10732A),.CK(CKA));
SDFF_X1 U_g1744A (.Q(g1744A),.SE(test_seA),.SI(g1209A),.D(g4239A),.CK(CKA));
SDFF_X1 U_g1558A (.Q(g1558A),.SE(test_seA),.SI(g1744A),.D(g6538A),.CK(CKA));
SDFF_X1 U_g695A (.Q(g695A),.SE(test_seA),.SI(g1558A),.D(g8887A),.CK(CKA));
SDFF_X1 U_g461A (.Q(g461A),.SE(test_seA),.SI(g695A),.D(g11372A),.CK(CKA));
SDFF_X1 U_g940A (.Q(g940A),.SE(test_seA),.SI(g461A),.D(g8260A),.CK(CKA));
SDFF_X1 U_g976A (.Q(g976A),.SE(test_seA),.SI(g940A),.D(g11391A),.CK(CKA));
SDFF_X1 U_g709A (.Q(g709A),.SE(test_seA),.SI(g976A),.D(g8432A),.CK(CKA));
SDFF_X1 U_g1092A (.Q(g1092A),.SE(test_seA),.SI(g709A),.D(g6088A),.CK(CKA));
SDFF_X1 U_g1574A (.Q(g1574A),.SE(test_seA),.SI(g1092A),.D(g6478A),.CK(CKA));
SDFF_X1 U_g1864A (.Q(g1864A),.SE(test_seA),.SI(g1574A),.D(g6795A),.CK(CKA));
SDFF_X1 U_g369A (.Q(g369A),.SE(test_seA),.SI(g1864A),.D(g11320A),.CK(CKA));
SDFF_X1 U_g1580A (.Q(g1580A),.SE(test_seA),.SI(g369A),.D(g6500A),.CK(CKA));
SDFF_X1 U_g1736A (.Q(g1736A),.SE(test_seA),.SI(g1580A),.D(g5392A),.CK(CKA));
SDFF_X1 U_g39A (.Q(g39A),.SE(test_seA),.SI(g1736A),.D(g10663A),.CK(CKA));
SDFF_X1 U_g1651A (.Q(g1651A),.SE(test_seA),.SI(g39A),.D(g10782A),.CK(CKA));
SDFF_X1 U_g1424A (.Q(g1424A),.SE(test_seA),.SI(g1651A),.D(g6216A),.CK(CKA));
SDFF_X1 U_g1737A (.Q(g1737A),.SE(test_seA),.SI(g1424A),.D(g1736A),.CK(CKA));
SDFF_X1 U_g1672A (.Q(g1672A),.SE(test_seA),.SI(g1737A),.D(g10858A),.CK(CKA));
SDFF_X1 U_g1077A (.Q(g1077A),.SE(test_seA),.SI(g1672A),.D(g5914A),.CK(CKA));
SDFF_X1 U_g1231A (.Q(g1231A),.SE(test_seA),.SI(g1077A),.D(g7590A),.CK(CKA));
SDFF_X1 U_g4A (.Q(g4A),.SE(test_seA),.SI(g1231A),.D(g6656A),.CK(CKA));
SDFF_X1 U_g774A (.Q(g774A),.SE(test_seA),.SI(g4A),.D(g6728A),.CK(CKA));
SDFF_X1 U_g1104A (.Q(g1104A),.SE(test_seA),.SI(g774A),.D(g5126A),.CK(CKA));
SDFF_X1 U_g1304A (.Q(g1304A),.SE(test_seA),.SI(g1104A),.D(g7290A),.CK(CKA));
SDFF_X1 U_g243A (.Q(g243A),.SE(test_seA),.SI(g1304A),.D(g6841A),.CK(CKA));
SDFF_X1 U_g1499A (.Q(g1499A),.SE(test_seA),.SI(g243A),.D(g8041A),.CK(CKA));
SDFF_X1 U_g1044A (.Q(g1044A),.SE(test_seA),.SI(g1499A),.D(g7106A),.CK(CKA));
SDFF_X1 U_g1444A (.Q(g1444A),.SE(test_seA),.SI(g1044A),.D(g8766A),.CK(CKA));
SDFF_X1 U_g757A (.Q(g757A),.SE(test_seA),.SI(g1444A),.D(g10788A),.CK(CKA));
SDFF_X1 U_g786A (.Q(g786A),.SE(test_seA),.SI(g757A),.D(g8019A),.CK(CKA));
SDFF_X1 U_g1543A (.Q(g1543A),.SE(test_seA),.SI(g786A),.D(g6545A),.CK(CKA));
SDFF_X1 U_g552A (.Q(g552A),.SE(test_seA),.SI(g1543A),.D(g10856A),.CK(CKA));
SDFF_X1 U_g315A (.Q(g315A),.SE(test_seA),.SI(g552A),.D(g256A),.CK(CKA));
SDFF_X1 U_g1534A (.Q(g1534A),.SE(test_seA),.SI(g315A),.D(g6533A),.CK(CKA));
SDFF_X1 U_g622A (.Q(g622A),.SE(test_seA),.SI(g1534A),.D(g8820A),.CK(CKA));
SDFF_X1 U_g1927A (.Q(g1927A),.SE(test_seA),.SI(g622A),.D(g8941A),.CK(CKA));
SDFF_X1 U_g1660A (.Q(g1660A),.SE(test_seA),.SI(g1927A),.D(g10859A),.CK(CKA));
SDFF_X1 U_g278A (.Q(g278A),.SE(test_seA),.SI(g1660A),.D(g6922A),.CK(CKA));
SDFF_X1 U_g1436A (.Q(g1436A),.SE(test_seA),.SI(g278A),.D(g8772A),.CK(CKA));
SDFF_X1 U_g718A (.Q(g718A),.SE(test_seA),.SI(g1436A),.D(g8433A),.CK(CKA));
SDFF_X1 U_g76A (.Q(g76A),.SE(test_seA),.SI(g718A),.D(g6526A),.CK(CKA));
SDFF_X1 U_g554A (.Q(g554A),.SE(test_seA),.SI(g76A),.D(g10793A),.CK(CKA));
SDFF_X1 U_g496A (.Q(g496A),.SE(test_seA),.SI(g554A),.D(g11333A),.CK(CKA));
SDFF_X1 U_g981A (.Q(g981A),.SE(test_seA),.SI(g496A),.D(g11392A),.CK(CKA));
SDFF_X1 U_g878A (.Q(g878A),.SE(test_seA),.SI(g981A),.D(g3506A),.CK(CKA));
SDFF_X1 U_g590A (.Q(g590A),.SE(test_seA),.SI(g878A),.D(g1713A),.CK(CKA));
SDFF_X1 U_g829A (.Q(g829A),.SE(test_seA),.SI(g590A),.D(g794A),.CK(CKA));
SDFF_X1 U_g1095A (.Q(g1095A),.SE(test_seA),.SI(g829A),.D(g6093A),.CK(CKA));
SDFF_X1 U_g704A (.Q(g704A),.SE(test_seA),.SI(g1095A),.D(g8889A),.CK(CKA));
SDFF_X1 U_g1265A (.Q(g1265A),.SE(test_seA),.SI(g704A),.D(g7302A),.CK(CKA));
SDFF_X1 U_g1786A (.Q(g1786A),.SE(test_seA),.SI(g1265A),.D(g6525A),.CK(CKA));
SDFF_X1 U_g682A (.Q(g682A),.SE(test_seA),.SI(g1786A),.D(g8429A),.CK(CKA));
SDFF_X1 U_g1296A (.Q(g1296A),.SE(test_seA),.SI(g682A),.D(g7292A),.CK(CKA));
SDFF_X1 U_g587A (.Q(g587A),.SE(test_seA),.SI(g1296A),.D(g104A),.CK(CKA));
SDFF_X1 U_g52A (.Q(g52A),.SE(test_seA),.SI(g587A),.D(g6621A),.CK(CKA));
SDFF_X1 U_g646A (.Q(g646A),.SE(test_seA),.SI(g52A),.D(g7134A),.CK(CKA));
SDFF_X1 U_g327A (.Q(g327A),.SE(test_seA),.SI(g646A),.D(g260A),.CK(CKA));
SDFF_X1 U_g1389A (.Q(g1389A),.SE(test_seA),.SI(g327A),.D(g6333A),.CK(CKA));
SDFF_X1 U_g1371A (.Q(g1371A),.SE(test_seA),.SI(g1389A),.D(g6826A),.CK(CKA));
SDFF_X1 U_g1956A (.Q(g1956A),.SE(test_seA),.SI(g1371A),.D(g1955A),.CK(CKA));
SDFF_X1 U_g1675A (.Q(g1675A),.SE(test_seA),.SI(g1956A),.D(g10860A),.CK(CKA));
SDFF_X1 U_g354A (.Q(g354A),.SE(test_seA),.SI(g1675A),.D(g11483A),.CK(CKA));
SDFF_X1 U_g113A (.Q(g113A),.SE(test_seA),.SI(g354A),.D(g6392A),.CK(CKA));
SDFF_X1 U_g639A (.Q(g639A),.SE(test_seA),.SI(g113A),.D(g7626A),.CK(CKA));
SDFF_X1 U_g1684A (.Q(g1684A),.SE(test_seA),.SI(g639A),.D(g10866A),.CK(CKA));
SDFF_X1 U_g1639A (.Q(g1639A),.SE(test_seA),.SI(g1684A),.D(g8193A),.CK(CKA));
SDFF_X1 U_g1791A (.Q(g1791A),.SE(test_seA),.SI(g1639A),.D(g6983A),.CK(CKA));
SDFF_X1 U_g248A (.Q(g248A),.SE(test_seA),.SI(g1791A),.D(g6839A),.CK(CKA));
SDFF_X1 U_g1707A (.Q(g1707A),.SE(test_seA),.SI(g248A),.D(g4076A),.CK(CKA));
SDFF_X1 U_g1759A (.Q(g1759A),.SE(test_seA),.SI(g1707A),.D(g4293A),.CK(CKA));
SDFF_X1 U_g351A (.Q(g351A),.SE(test_seA),.SI(g1759A),.D(g11482A),.CK(CKA));
SDFF_X1 U_g1957A (.Q(g1957A),.SE(test_seA),.SI(g351A),.D(g1956A),.CK(CKA));
SDFF_X1 U_g1604A (.Q(g1604A),.SE(test_seA),.SI(g1957A),.D(g6507A),.CK(CKA));
SDFF_X1 U_g1098A (.Q(g1098A),.SE(test_seA),.SI(g1604A),.D(g6096A),.CK(CKA));
SDFF_X1 U_g932A (.Q(g932A),.SE(test_seA),.SI(g1098A),.D(g8250A),.CK(CKA));
SDFF_X1 U_g126A (.Q(g126A),.SE(test_seA),.SI(g932A),.D(I8503A),.CK(CKA));
SDFF_X1 U_g1896A (.Q(g1896A),.SE(test_seA),.SI(g126A),.D(g8282A),.CK(CKA));
SDFF_X1 U_g736A (.Q(g736A),.SE(test_seA),.SI(g1896A),.D(g8435A),.CK(CKA));
SDFF_X1 U_g1019A (.Q(g1019A),.SE(test_seA),.SI(g736A),.D(g6924A),.CK(CKA));
SDFF_X1 U_g1362A (.Q(g1362A),.SE(test_seA),.SI(g1019A),.D(g6819A),.CK(CKA));
SDFF_X1 U_g745A (.Q(g745A),.SE(test_seA),.SI(g1362A),.D(g746A),.CK(CKA));
SDFF_X1 U_g1419A (.Q(g1419A),.SE(test_seA),.SI(g745A),.D(g6244A),.CK(CKA));
SDFF_X1 U_g58A (.Q(g58A),.SE(test_seA),.SI(g1419A),.D(g6627A),.CK(CKA));
SDFF_X1 U_g32A (.Q(g32A),.SE(test_seA),.SI(g58A),.D(g11286A),.CK(CKA));
SDFF_X1 U_g876A (.Q(g876A),.SE(test_seA),.SI(g32A),.D(g878A),.CK(CKA));
SDFF_X1 U_g1086A (.Q(g1086A),.SE(test_seA),.SI(g876A),.D(g6071A),.CK(CKA));
SDFF_X1 U_g1486A (.Q(g1486A),.SE(test_seA),.SI(g1086A),.D(g8046A),.CK(CKA));
SDFF_X1 U_g1730A (.Q(g1730A),.SE(test_seA),.SI(g1486A),.D(g10707A),.CK(CKA));
SDFF_X1 U_g1504A (.Q(g1504A),.SE(test_seA),.SI(g1730A),.D(g6198A),.CK(CKA));
SDFF_X1 U_g1470A (.Q(g1470A),.SE(test_seA),.SI(g1504A),.D(g8051A),.CK(CKA));
SDFF_X1 U_g822A (.Q(g822A),.SE(test_seA),.SI(g1470A),.D(g8024A),.CK(CKA));
SDFF_X1 U_g583A (.Q(g583A),.SE(test_seA),.SI(g822A),.D(g29A),.CK(CKA));
SDFF_X1 U_g1678A (.Q(g1678A),.SE(test_seA),.SI(g583A),.D(g10862A),.CK(CKA));
SDFF_X1 U_g174A (.Q(g174A),.SE(test_seA),.SI(g1678A),.D(g8050A),.CK(CKA));
SDFF_X1 U_g1766A (.Q(g1766A),.SE(test_seA),.SI(g174A),.D(g7133A),.CK(CKA));
SDFF_X1 U_g1801A (.Q(g1801A),.SE(test_seA),.SI(g1766A),.D(g7930A),.CK(CKA));
SDFF_X1 U_g186A (.Q(g186A),.SE(test_seA),.SI(g1801A),.D(g6832A),.CK(CKA));
SDFF_X1 U_g959A (.Q(g959A),.SE(test_seA),.SI(g186A),.D(g11308A),.CK(CKA));
SDFF_X1 U_g1169A (.Q(g1169A),.SE(test_seA),.SI(g959A),.D(g5189A),.CK(CKA));
SDFF_X1 U_g1007A (.Q(g1007A),.SE(test_seA),.SI(g1169A),.D(g6918A),.CK(CKA));
SDFF_X1 U_g1407A (.Q(g1407A),.SE(test_seA),.SI(g1007A),.D(g8769A),.CK(CKA));
SDFF_X1 U_g1059A (.Q(g1059A),.SE(test_seA),.SI(g1407A),.D(g7236A),.CK(CKA));
SDFF_X1 U_g1868A (.Q(g1868A),.SE(test_seA),.SI(g1059A),.D(g6909A),.CK(CKA));
SDFF_X1 U_g758A (.Q(g758A),.SE(test_seA),.SI(g1868A),.D(g4940A),.CK(CKA));
SDFF_X1 U_g1718A (.Q(g1718A),.SE(test_seA),.SI(g758A),.D(g5404A),.CK(CKA));
SDFF_X1 U_g396A (.Q(g396A),.SE(test_seA),.SI(g1718A),.D(g11265A),.CK(CKA));
SDFF_X1 U_g1015A (.Q(g1015A),.SE(test_seA),.SI(g396A),.D(g6930A),.CK(CKA));
SDFF_X1 U_g38A (.Q(g38A),.SE(test_seA),.SI(g1015A),.D(g10726A),.CK(CKA));
SDFF_X1 U_g632A (.Q(g632A),.SE(test_seA),.SI(g38A),.D(g4891A),.CK(CKA));
SDFF_X1 U_g1415A (.Q(g1415A),.SE(test_seA),.SI(g632A),.D(g6224A),.CK(CKA));
SDFF_X1 U_g1227A (.Q(g1227A),.SE(test_seA),.SI(g1415A),.D(g7586A),.CK(CKA));
SDFF_X1 U_g1721A (.Q(g1721A),.SE(test_seA),.SI(g1227A),.D(g10770A),.CK(CKA));
SDFF_X1 U_g882A (.Q(g882A),.SE(test_seA),.SI(g1721A),.D(g883A),.CK(CKA));
SDFF_X1 U_g16A (.Q(g16A),.SE(test_seA),.SI(g882A),.D(g3524A),.CK(CKA));
SDFF_X1 U_g284A (.Q(g284A),.SE(test_seA),.SI(g16A),.D(g6934A),.CK(CKA));
SDFF_X1 U_g426A (.Q(g426A),.SE(test_seA),.SI(g284A),.D(g11256A),.CK(CKA));
SDFF_X1 U_g219A (.Q(g219A),.SE(test_seA),.SI(g426A),.D(g6824A),.CK(CKA));
SDFF_X1 U_g1216A (.Q(g1216A),.SE(test_seA),.SI(g219A),.D(g1360A),.CK(CKA));
SDFF_X1 U_g806A (.Q(g806A),.SE(test_seA),.SI(g1216A),.D(g6126A),.CK(CKA));
SDFF_X1 U_g1428A (.Q(g1428A),.SE(test_seA),.SI(g806A),.D(g8767A),.CK(CKA));
SDFF_X1 U_g579A (.Q(g579A),.SE(test_seA),.SI(g1428A),.D(g102A),.CK(CKA));
SDFF_X1 U_g1564A (.Q(g1564A),.SE(test_seA),.SI(g579A),.D(g6546A),.CK(CKA));
SDFF_X1 U_g1741A (.Q(g1741A),.SE(test_seA),.SI(g1564A),.D(g4238A),.CK(CKA));
SDFF_X1 U_g225A (.Q(g225A),.SE(test_seA),.SI(g1741A),.D(g6823A),.CK(CKA));
SDFF_X1 U_g281A (.Q(g281A),.SE(test_seA),.SI(g225A),.D(g6928A),.CK(CKA));
SDFF_X1 U_g1308A (.Q(g1308A),.SE(test_seA),.SI(g281A),.D(g11602A),.CK(CKA));
SDFF_X1 U_g611A (.Q(g611A),.SE(test_seA),.SI(g1308A),.D(g9721A),.CK(CKA));
SDFF_X1 U_g631A (.Q(g631A),.SE(test_seA),.SI(g611A),.D(g4890A),.CK(CKA));
SDFF_X1 U_g1217A (.Q(g1217A),.SE(test_seA),.SI(g631A),.D(g9525A),.CK(CKA));
SDFF_X1 U_g1589A (.Q(g1589A),.SE(test_seA),.SI(g1217A),.D(g6524A),.CK(CKA));
SDFF_X1 U_g1466A (.Q(g1466A),.SE(test_seA),.SI(g1589A),.D(g8045A),.CK(CKA));
SDFF_X1 U_g1571A (.Q(g1571A),.SE(test_seA),.SI(g1466A),.D(g6469A),.CK(CKA));
SDFF_X1 U_g1861A (.Q(g1861A),.SE(test_seA),.SI(g1571A),.D(g6471A),.CK(CKA));
SDFF_X1 U_g1365A (.Q(g1365A),.SE(test_seA),.SI(g1861A),.D(g6821A),.CK(CKA));
SDFF_X1 U_g1448A (.Q(g1448A),.SE(test_seA),.SI(g1365A),.D(g11514A),.CK(CKA));
SDFF_X1 U_g1711A (.Q(g1711A),.SE(test_seA),.SI(g1448A),.D(g5403A),.CK(CKA));
SDFF_X1 U_g1133A (.Q(g1133A),.SE(test_seA),.SI(g1711A),.D(g4480A),.CK(CKA));
SDFF_X1 U_g1333A (.Q(g1333A),.SE(test_seA),.SI(g1133A),.D(g11610A),.CK(CKA));
SDFF_X1 U_g153A (.Q(g153A),.SE(test_seA),.SI(g1333A),.D(g7843A),.CK(CKA));
SDFF_X1 U_g962A (.Q(g962A),.SE(test_seA),.SI(g153A),.D(g11310A),.CK(CKA));
SDFF_X1 U_g766A (.Q(g766A),.SE(test_seA),.SI(g962A),.D(g5536A),.CK(CKA));
SDFF_X1 U_g588A (.Q(g588A),.SE(test_seA),.SI(g766A),.D(g28A),.CK(CKA));
SDFF_X1 U_g486A (.Q(g486A),.SE(test_seA),.SI(g588A),.D(g11331A),.CK(CKA));
SDFF_X1 U_g471A (.Q(g471A),.SE(test_seA),.SI(g486A),.D(g11380A),.CK(CKA));
SDFF_X1 U_g1397A (.Q(g1397A),.SE(test_seA),.SI(g471A),.D(g6838A),.CK(CKA));
SDFF_X1 U_g580A (.Q(g580A),.SE(test_seA),.SI(g1397A),.D(g103A),.CK(CKA));
SDFF_X1 U_g1950A (.Q(g1950A),.SE(test_seA),.SI(g580A),.D(g8288A),.CK(CKA));
SDFF_X1 U_g756A (.Q(g756A),.SE(test_seA),.SI(g1950A),.D(g755A),.CK(CKA));
SDFF_X1 U_g635A (.Q(g635A),.SE(test_seA),.SI(g756A),.D(g4892A),.CK(CKA));
SDFF_X1 U_g1101A (.Q(g1101A),.SE(test_seA),.SI(g635A),.D(g5390A),.CK(CKA));
SDFF_X1 U_g549A (.Q(g549A),.SE(test_seA),.SI(g1101A),.D(g10855A),.CK(CKA));
SDFF_X1 U_g1041A (.Q(g1041A),.SE(test_seA),.SI(g549A),.D(g7258A),.CK(CKA));
SDFF_X1 U_g105A (.Q(g105A),.SE(test_seA),.SI(g1041A),.D(g10898A),.CK(CKA));
SDFF_X1 U_g1669A (.Q(g1669A),.SE(test_seA),.SI(g105A),.D(g10865A),.CK(CKA));
SDFF_X1 U_g1368A (.Q(g1368A),.SE(test_seA),.SI(g1669A),.D(g6822A),.CK(CKA));
SDFF_X1 U_g1531A (.Q(g1531A),.SE(test_seA),.SI(g1368A),.D(g6528A),.CK(CKA));
SDFF_X1 U_g1458A (.Q(g1458A),.SE(test_seA),.SI(g1531A),.D(g6180A),.CK(CKA));
SDFF_X1 U_g572A (.Q(g572A),.SE(test_seA),.SI(g1458A),.D(g10718A),.CK(CKA));
SDFF_X1 U_g1011A (.Q(g1011A),.SE(test_seA),.SI(g572A),.D(g6912A),.CK(CKA));
SDFF_X1 U_g33A (.Q(g33A),.SE(test_seA),.SI(g1011A),.D(g10719A),.CK(CKA));
SDFF_X1 U_g1411A (.Q(g1411A),.SE(test_seA),.SI(g33A),.D(g6234A),.CK(CKA));
SDFF_X1 U_g1074A (.Q(g1074A),.SE(test_seA),.SI(g1411A),.D(g6099A),.CK(CKA));
SDFF_X1 U_g444A (.Q(g444A),.SE(test_seA),.SI(g1074A),.D(g11259A),.CK(CKA));
SDFF_X1 U_g1474A (.Q(g1474A),.SE(test_seA),.SI(g444A),.D(g8039A),.CK(CKA));
SDFF_X1 U_g1080A (.Q(g1080A),.SE(test_seA),.SI(g1474A),.D(g6059A),.CK(CKA));
SDFF_X1 U_g1713A (.Q(g1713A),.SE(test_seA),.SI(g1080A),.D(g5396A),.CK(CKA));
SDFF_X1 U_g333A (.Q(g333A),.SE(test_seA),.SI(g1713A),.D(g262A),.CK(CKA));
SDFF_X1 U_g269A (.Q(g269A),.SE(test_seA),.SI(g333A),.D(g6906A),.CK(CKA));
SDFF_X1 U_g401A (.Q(g401A),.SE(test_seA),.SI(g269A),.D(g11266A),.CK(CKA));
SDFF_X1 U_g1857A (.Q(g1857A),.SE(test_seA),.SI(g401A),.D(g11294A),.CK(CKA));
SDFF_X1 U_g9A (.Q(g9A),.SE(test_seA),.SI(g1857A),.D(g5421A),.CK(CKA));
SDFF_X1 U_g664A (.Q(g664A),.SE(test_seA),.SI(g9A),.D(g8649A),.CK(CKA));
SDFF_X1 U_g965A (.Q(g965A),.SE(test_seA),.SI(g664A),.D(g11312A),.CK(CKA));
SDFF_X1 U_g1400A (.Q(g1400A),.SE(test_seA),.SI(g965A),.D(g6840A),.CK(CKA));
SDFF_X1 U_g309A (.Q(g309A),.SE(test_seA),.SI(g1400A),.D(g254A),.CK(CKA));
SDFF_X1 U_g814A (.Q(g814A),.SE(test_seA),.SI(g309A),.D(g7202A),.CK(CKA));
SDFF_X1 U_g231A (.Q(g231A),.SE(test_seA),.SI(g814A),.D(g6834A),.CK(CKA));
SDFF_X1 U_g557A (.Q(g557A),.SE(test_seA),.SI(g231A),.D(g10795A),.CK(CKA));
SDFF_X1 U_g586A (.Q(g586A),.SE(test_seA),.SI(g557A),.D(g103A),.CK(CKA));
SDFF_X1 U_g869A (.Q(g869A),.SE(test_seA),.SI(g586A),.D(g875A),.CK(CKA));
SDFF_X1 U_g1383A (.Q(g1383A),.SE(test_seA),.SI(g869A),.D(g6831A),.CK(CKA));
SDFF_X1 U_g158A (.Q(g158A),.SE(test_seA),.SI(g1383A),.D(g8060A),.CK(CKA));
SDFF_X1 U_g627A (.Q(g627A),.SE(test_seA),.SI(g158A),.D(g4893A),.CK(CKA));
SDFF_X1 U_g1023A (.Q(g1023A),.SE(test_seA),.SI(g627A),.D(g7244A),.CK(CKA));
SDFF_X1 U_g259A (.Q(g259A),.SE(test_seA),.SI(g1023A),.D(g6026A),.CK(CKA));
SDFF_X1 U_g1361A (.Q(g1361A),.SE(test_seA),.SI(g259A),.D(g1206A),.CK(CKA));
SDFF_X1 U_g1327A (.Q(g1327A),.SE(test_seA),.SI(g1361A),.D(g11608A),.CK(CKA));
SDFF_X1 U_g654A (.Q(g654A),.SE(test_seA),.SI(g1327A),.D(g7660A),.CK(CKA));
SDFF_X1 U_g293A (.Q(g293A),.SE(test_seA),.SI(g654A),.D(g6911A),.CK(CKA));
SDFF_X1 U_g1346A (.Q(g1346A),.SE(test_seA),.SI(g293A),.D(g11640A),.CK(CKA));
SDFF_X1 U_g1633A (.Q(g1633A),.SE(test_seA),.SI(g1346A),.D(g8777A),.CK(CKA));
SDFF_X1 U_g1753A (.Q(g1753A),.SE(test_seA),.SI(g1633A),.D(g4274A),.CK(CKA));
SDFF_X1 U_g1508A (.Q(g1508A),.SE(test_seA),.SI(g1753A),.D(g6215A),.CK(CKA));
SDFF_X1 U_g1240A (.Q(g1240A),.SE(test_seA),.SI(g1508A),.D(g7297A),.CK(CKA));
SDFF_X1 U_g538A (.Q(g538A),.SE(test_seA),.SI(g1240A),.D(g11326A),.CK(CKA));
SDFF_X1 U_g416A (.Q(g416A),.SE(test_seA),.SI(g538A),.D(g11269A),.CK(CKA));
SDFF_X1 U_g542A (.Q(g542A),.SE(test_seA),.SI(g416A),.D(g11325A),.CK(CKA));
SDFF_X1 U_g1681A (.Q(g1681A),.SE(test_seA),.SI(g542A),.D(g10864A),.CK(CKA));
SDFF_X1 U_g374A (.Q(g374A),.SE(test_seA),.SI(g1681A),.D(g11290A),.CK(CKA));
SDFF_X1 U_g563A (.Q(g563A),.SE(test_seA),.SI(g374A),.D(g10798A),.CK(CKA));
SDFF_X1 U_g1914A (.Q(g1914A),.SE(test_seA),.SI(g563A),.D(g8284A),.CK(CKA));
SDFF_X1 U_g530A (.Q(g530A),.SE(test_seA),.SI(g1914A),.D(g11328A),.CK(CKA));
SDFF_X1 U_g575A (.Q(g575A),.SE(test_seA),.SI(g530A),.D(g10800A),.CK(CKA));
SDFF_X1 U_g1936A (.Q(g1936A),.SE(test_seA),.SI(g575A),.D(g8944A),.CK(CKA));
SDFF_X1 U_g55A (.Q(g55A),.SE(test_seA),.SI(g1936A),.D(g7183A),.CK(CKA));
SDFF_X1 U_g1117A (.Q(g1117A),.SE(test_seA),.SI(g55A),.D(g4465A),.CK(CKA));
SDFF_X1 U_g1317A (.Q(g1317A),.SE(test_seA),.SI(g1117A),.D(g1356A),.CK(CKA));
SDFF_X1 U_g357A (.Q(g357A),.SE(test_seA),.SI(g1317A),.D(g11484A),.CK(CKA));
SDFF_X1 U_g386A (.Q(g386A),.SE(test_seA),.SI(g357A),.D(g11263A),.CK(CKA));
SDFF_X1 U_g1601A (.Q(g1601A),.SE(test_seA),.SI(g386A),.D(g6501A),.CK(CKA));
SDFF_X1 U_g553A (.Q(g553A),.SE(test_seA),.SI(g1601A),.D(g10857A),.CK(CKA));
SDFF_X1 U_g166A (.Q(g166A),.SE(test_seA),.SI(g553A),.D(g6757A),.CK(CKA));
SDFF_X1 U_g501A (.Q(g501A),.SE(test_seA),.SI(g166A),.D(g11334A),.CK(CKA));
SDFF_X1 U_g262A (.Q(g262A),.SE(test_seA),.SI(g501A),.D(g6042A),.CK(CKA));
SDFF_X1 U_g1840A (.Q(g1840A),.SE(test_seA),.SI(g262A),.D(g8384A),.CK(CKA));
SDFF_X1 U_g70A (.Q(g70A),.SE(test_seA),.SI(g1840A),.D(g6653A),.CK(CKA));
SDFF_X1 U_g318A (.Q(g318A),.SE(test_seA),.SI(g70A),.D(g257A),.CK(CKA));
SDFF_X1 U_g1356A (.Q(g1356A),.SE(test_seA),.SI(g318A),.D(g5763A),.CK(CKA));
SDFF_X1 U_g794A (.Q(g794A),.SE(test_seA),.SI(g1356A),.D(g5849A),.CK(CKA));
SDFF_X1 U_g36A (.Q(g36A),.SE(test_seA),.SI(g794A),.D(g10722A),.CK(CKA));
SDFF_X1 U_g302A (.Q(g302A),.SE(test_seA),.SI(g36A),.D(g6929A),.CK(CKA));
SDFF_X1 U_g342A (.Q(g342A),.SE(test_seA),.SI(g302A),.D(g11488A),.CK(CKA));
SDFF_X1 U_g1250A (.Q(g1250A),.SE(test_seA),.SI(g342A),.D(g7299A),.CK(CKA));
SDFF_X1 U_g1163A (.Q(g1163A),.SE(test_seA),.SI(g1250A),.D(g4330A),.CK(CKA));
SDFF_X1 U_g1810A (.Q(g1810A),.SE(test_seA),.SI(g1163A),.D(g1958A),.CK(CKA));
SDFF_X1 U_g1032A (.Q(g1032A),.SE(test_seA),.SI(g1810A),.D(g7257A),.CK(CKA));
SDFF_X1 U_g1432A (.Q(g1432A),.SE(test_seA),.SI(g1032A),.D(g8775A),.CK(CKA));
SDFF_X1 U_g1053A (.Q(g1053A),.SE(test_seA),.SI(g1432A),.D(g7225A),.CK(CKA));
SDFF_X1 U_g1453A (.Q(g1453A),.SE(test_seA),.SI(g1053A),.D(g5770A),.CK(CKA));
SDFF_X1 U_g363A (.Q(g363A),.SE(test_seA),.SI(g1453A),.D(g11486A),.CK(CKA));
SDFF_X1 U_g330A (.Q(g330A),.SE(test_seA),.SI(g363A),.D(g261A),.CK(CKA));
SDFF_X1 U_g1157A (.Q(g1157A),.SE(test_seA),.SI(g330A),.D(g4338A),.CK(CKA));
SDFF_X1 U_g1357A (.Q(g1357A),.SE(test_seA),.SI(g1157A),.D(g4500A),.CK(CKA));
SDFF_X1 U_g35A (.Q(g35A),.SE(test_seA),.SI(g1357A),.D(g10721A),.CK(CKA));
SDFF_X1 U_g928A (.Q(g928A),.SE(test_seA),.SI(g35A),.D(g8147A),.CK(CKA));
SDFF_X1 U_g261A (.Q(g261A),.SE(test_seA),.SI(g928A),.D(g6038A),.CK(CKA));
SDFF_X1 U_g516A (.Q(g516A),.SE(test_seA),.SI(g261A),.D(g11337A),.CK(CKA));
SDFF_X1 U_g254A (.Q(g254A),.SE(test_seA),.SI(g516A),.D(g6045A),.CK(CKA));
SDFF_X1 U_g778A (.Q(g778A),.SE(test_seA),.SI(g254A),.D(g7191A),.CK(CKA));
SDFF_X1 U_g861A (.Q(g861A),.SE(test_seA),.SI(g778A),.D(g826A),.CK(CKA));
SDFF_X1 U_g1627A (.Q(g1627A),.SE(test_seA),.SI(g861A),.D(g8774A),.CK(CKA));
SDFF_X1 U_g1292A (.Q(g1292A),.SE(test_seA),.SI(g1627A),.D(g7293A),.CK(CKA));
SDFF_X1 U_g290A (.Q(g290A),.SE(test_seA),.SI(g1292A),.D(g6907A),.CK(CKA));
SDFF_X1 U_g1850A (.Q(g1850A),.SE(test_seA),.SI(g290A),.D(g4903A),.CK(CKA));
SDFF_X1 U_g770A (.Q(g770A),.SE(test_seA),.SI(g1850A),.D(g6123A),.CK(CKA));
SDFF_X1 U_g1583A (.Q(g1583A),.SE(test_seA),.SI(g770A),.D(g6506A),.CK(CKA));
SDFF_X1 U_g466A (.Q(g466A),.SE(test_seA),.SI(g1583A),.D(g11376A),.CK(CKA));
SDFF_X1 U_g1561A (.Q(g1561A),.SE(test_seA),.SI(g466A),.D(g6542A),.CK(CKA));
SDFF_X1 U_g1527A (.Q(g1527A),.SE(test_seA),.SI(g1561A),.D(I8503A),.CK(CKA));
SDFF_X1 U_g1546A (.Q(g1546A),.SE(test_seA),.SI(g1527A),.D(g6551A),.CK(CKA));
SDFF_X1 U_g287A (.Q(g287A),.SE(test_seA),.SI(g1546A),.D(g6901A),.CK(CKA));
SDFF_X1 U_g560A (.Q(g560A),.SE(test_seA),.SI(g287A),.D(g10797A),.CK(CKA));
SDFF_X1 U_g617A (.Q(g617A),.SE(test_seA),.SI(g560A),.D(g8505A),.CK(CKA));
SDFF_X1 U_g17A (.Q(g17A),.SE(test_seA),.SI(g617A),.D(g4117A),.CK(CKA));
SDFF_X1 U_g336A (.Q(g336A),.SE(test_seA),.SI(g17A),.D(g11647A),.CK(CKA));
SDFF_X1 U_g456A (.Q(g456A),.SE(test_seA),.SI(g336A),.D(g11340A),.CK(CKA));
SDFF_X1 U_g305A (.Q(g305A),.SE(test_seA),.SI(g456A),.D(g253A),.CK(CKA));
SDFF_X1 U_g345A (.Q(g345A),.SE(test_seA),.SI(g305A),.D(g11625A),.CK(CKA));
SDFF_X1 U_g8A (.Q(g8A),.SE(test_seA),.SI(g345A),.D(g636A),.CK(CKA));
SDFF_X1 U_g1771A (.Q(g1771A),.SE(test_seA),.SI(g8A),.D(g6502A),.CK(CKA));
SDFF_X1 U_g865A (.Q(g865A),.SE(test_seA),.SI(g1771A),.D(g7981A),.CK(CKA));
SDFF_X1 U_g255A (.Q(g255A),.SE(test_seA),.SI(g865A),.D(g6049A),.CK(CKA));
SDFF_X1 U_g1945A (.Q(g1945A),.SE(test_seA),.SI(g255A),.D(g8945A),.CK(CKA));
SDFF_X1 U_g1738A (.Q(g1738A),.SE(test_seA),.SI(g1945A),.D(g4231A),.CK(CKA));
SDFF_X1 U_g1478A (.Q(g1478A),.SE(test_seA),.SI(g1738A),.D(g8040A),.CK(CKA));
SDFF_X1 U_g1035A (.Q(g1035A),.SE(test_seA),.SI(g1478A),.D(g7203A),.CK(CKA));
SDFF_X1 U_g1959A (.Q(g1959A),.SE(test_seA),.SI(g1035A),.D(I5254A),.CK(CKA));
SDFF_X1 U_g1690A (.Q(g1690A),.SE(test_seA),.SI(g1959A),.D(g6155A),.CK(CKA));
SDFF_X1 U_g1482A (.Q(g1482A),.SE(test_seA),.SI(g1690A),.D(g8043A),.CK(CKA));
SDFF_X1 U_g1110A (.Q(g1110A),.SE(test_seA),.SI(g1482A),.D(g5173A),.CK(CKA));
SDFF_X1 U_g296A (.Q(g296A),.SE(test_seA),.SI(g1110A),.D(g6916A),.CK(CKA));
SDFF_X1 U_g1663A (.Q(g1663A),.SE(test_seA),.SI(g296A),.D(g10861A),.CK(CKA));
SDFF_X1 U_g700A (.Q(g700A),.SE(test_seA),.SI(g1663A),.D(g8431A),.CK(CKA));
SDFF_X1 U_g1762A (.Q(g1762A),.SE(test_seA),.SI(g700A),.D(g4309A),.CK(CKA));
SDFF_X1 U_g360A (.Q(g360A),.SE(test_seA),.SI(g1762A),.D(g11485A),.CK(CKA));
SDFF_X1 U_g192A (.Q(g192A),.SE(test_seA),.SI(g360A),.D(g6334A),.CK(CKA));
SDFF_X1 U_g1657A (.Q(g1657A),.SE(test_seA),.SI(g192A),.D(g10767A),.CK(CKA));
SDFF_X1 U_g722A (.Q(g722A),.SE(test_seA),.SI(g1657A),.D(g8923A),.CK(CKA));
SDFF_X1 U_g61A (.Q(g61A),.SE(test_seA),.SI(g722A),.D(g7189A),.CK(CKA));
SDFF_X1 U_g566A (.Q(g566A),.SE(test_seA),.SI(g61A),.D(g10799A),.CK(CKA));
SDFF_X1 U_g1394A (.Q(g1394A),.SE(test_seA),.SI(g566A),.D(g6747A),.CK(CKA));
SDFF_X1 U_g1089A (.Q(g1089A),.SE(test_seA),.SI(g1394A),.D(g6080A),.CK(CKA));
SDFF_X1 U_g883A (.Q(g883A),.SE(test_seA),.SI(g1089A),.D(g3381A),.CK(CKA));
SDFF_X1 U_g1071A (.Q(g1071A),.SE(test_seA),.SI(g883A),.D(g5910A),.CK(CKA));
SDFF_X1 U_g986A (.Q(g986A),.SE(test_seA),.SI(g1071A),.D(g11393A),.CK(CKA));
SDFF_X1 U_g971A (.Q(g971A),.SE(test_seA),.SI(g986A),.D(g11349A),.CK(CKA));
SDFF_X1 U_g1955A (.Q(g1955A),.SE(test_seA),.SI(g971A),.D(g83A),.CK(CKA));
SDFF_X1 U_g143A (.Q(g143A),.SE(test_seA),.SI(g1955A),.D(g6439A),.CK(CKA));
SDFF_X1 U_g1814A (.Q(g1814A),.SE(test_seA),.SI(g143A),.D(g9266A),.CK(CKA));
SDFF_X1 U_g1038A (.Q(g1038A),.SE(test_seA),.SI(g1814A),.D(g7245A),.CK(CKA));
SDFF_X1 U_g1212A (.Q(g1212A),.SE(test_seA),.SI(g1038A),.D(g1217A),.CK(CKA));
SDFF_X1 U_g1918A (.Q(g1918A),.SE(test_seA),.SI(g1212A),.D(g8940A),.CK(CKA));
SDFF_X1 U_g782A (.Q(g782A),.SE(test_seA),.SI(g1918A),.D(g7705A),.CK(CKA));
SDFF_X1 U_g1822A (.Q(g1822A),.SE(test_seA),.SI(g782A),.D(g9269A),.CK(CKA));
SDFF_X1 U_g237A (.Q(g237A),.SE(test_seA),.SI(g1822A),.D(g6820A),.CK(CKA));
SDFF_X1 U_g746A (.Q(g746A),.SE(test_seA),.SI(g237A),.D(g756A),.CK(CKA));
SDFF_X1 U_g1062A (.Q(g1062A),.SE(test_seA),.SI(g746A),.D(g7240A),.CK(CKA));
SDFF_X1 U_g1462A (.Q(g1462A),.SE(test_seA),.SI(g1062A),.D(g8042A),.CK(CKA));
SDFF_X1 U_g178A (.Q(g178A),.SE(test_seA),.SI(g1462A),.D(g6759A),.CK(CKA));
SDFF_X1 U_g366A (.Q(g366A),.SE(test_seA),.SI(g178A),.D(g11487A),.CK(CKA));
SDFF_X1 U_g837A (.Q(g837A),.SE(test_seA),.SI(g366A),.D(g802A),.CK(CKA));
SDFF_X1 U_g599A (.Q(g599A),.SE(test_seA),.SI(g837A),.D(g9124A),.CK(CKA));
SDFF_X1 U_g1854A (.Q(g1854A),.SE(test_seA),.SI(g599A),.D(g11293A),.CK(CKA));
SDFF_X1 U_g944A (.Q(g944A),.SE(test_seA),.SI(g1854A),.D(g11298A),.CK(CKA));
SDFF_X1 U_g1941A (.Q(g1941A),.SE(test_seA),.SI(g944A),.D(g8287A),.CK(CKA));
SDFF_X1 U_g170A (.Q(g170A),.SE(test_seA),.SI(g1941A),.D(g8047A),.CK(CKA));
SDFF_X1 U_g1520A (.Q(g1520A),.SE(test_seA),.SI(g170A),.D(g6205A),.CK(CKA));
SDFF_X1 U_g686A (.Q(g686A),.SE(test_seA),.SI(g1520A),.D(g8885A),.CK(CKA));
SDFF_X1 U_g953A (.Q(g953A),.SE(test_seA),.SI(g686A),.D(g11305A),.CK(CKA));
SDFF_X1 U_g1958A (.Q(g1958A),.SE(test_seA),.SI(g953A),.D(g5556A),.CK(CKA));
SDFF_X1 U_g40A (.Q(g40A),.SE(test_seA),.SI(g1958A),.D(g10664A),.CK(CKA));
SDFF_X1 U_g1765A (.Q(g1765A),.SE(test_seA),.SI(g40A),.D(g2478A),.CK(CKA));
SDFF_X1 U_g1733A (.Q(g1733A),.SE(test_seA),.SI(g1765A),.D(g10711A),.CK(CKA));
SDFF_X1 U_g1270A (.Q(g1270A),.SE(test_seA),.SI(g1733A),.D(g7303A),.CK(CKA));
SDFF_X1 U_g1610A (.Q(g1610A),.SE(test_seA),.SI(g1270A),.D(g5194A),.CK(CKA));
SDFF_X1 U_g1796A (.Q(g1796A),.SE(test_seA),.SI(g1610A),.D(g7541A),.CK(CKA));
SDFF_X1 U_g1324A (.Q(g1324A),.SE(test_seA),.SI(g1796A),.D(g11607A),.CK(CKA));
SDFF_X1 U_g1540A (.Q(g1540A),.SE(test_seA),.SI(g1324A),.D(g6541A),.CK(CKA));
SDFF_X1 U_g1377A (.Q(g1377A),.SE(test_seA),.SI(g1540A),.D(g6827A),.CK(CKA));
SDFF_X1 U_g1206A (.Q(g1206A),.SE(test_seA),.SI(g1377A),.D(g4114A),.CK(CKA));
SDFF_X1 U_g491A (.Q(g491A),.SE(test_seA),.SI(g1206A),.D(g11332A),.CK(CKA));
SDFF_X1 U_g1849A (.Q(g1849A),.SE(test_seA),.SI(g491A),.D(g4902A),.CK(CKA));
SDFF_X1 U_g213A (.Q(g213A),.SE(test_seA),.SI(g1849A),.D(g6828A),.CK(CKA));
SDFF_X1 U_g1781A (.Q(g1781A),.SE(test_seA),.SI(g213A),.D(g6516A),.CK(CKA));
SDFF_X1 U_g1900A (.Q(g1900A),.SE(test_seA),.SI(g1781A),.D(g8938A),.CK(CKA));
SDFF_X1 U_g1245A (.Q(g1245A),.SE(test_seA),.SI(g1900A),.D(g7298A),.CK(CKA));
SDFF_X1 U_g108A (.Q(g108A),.SE(test_seA),.SI(g1245A),.D(g11561A),.CK(CKA));
SDFF_X1 U_g630A (.Q(g630A),.SE(test_seA),.SI(g108A),.D(g6672A),.CK(CKA));
SDFF_X1 U_g148A (.Q(g148A),.SE(test_seA),.SI(g630A),.D(g8048A),.CK(CKA));
SDFF_X1 U_g833A (.Q(g833A),.SE(test_seA),.SI(g148A),.D(g798A),.CK(CKA));
SDFF_X1 U_g1923A (.Q(g1923A),.SE(test_seA),.SI(g833A),.D(g8285A),.CK(CKA));
SDFF_X1 U_g936A (.Q(g936A),.SE(test_seA),.SI(g1923A),.D(g8254A),.CK(CKA));
SDFF_X1 U_g1215A (.Q(g1215A),.SE(test_seA),.SI(g936A),.D(g5229A),.CK(CKA));
SDFF_X1 U_g1314A (.Q(g1314A),.SE(test_seA),.SI(g1215A),.D(g11604A),.CK(CKA));
SDFF_X1 U_g849A (.Q(g849A),.SE(test_seA),.SI(g1314A),.D(g814A),.CK(CKA));
SDFF_X1 U_g1336A (.Q(g1336A),.SE(test_seA),.SI(g849A),.D(g11636A),.CK(CKA));
SDFF_X1 U_g272A (.Q(g272A),.SE(test_seA),.SI(g1336A),.D(g6910A),.CK(CKA));
SDFF_X1 U_g1806A (.Q(g1806A),.SE(test_seA),.SI(g272A),.D(g8173A),.CK(CKA));
SDFF_X1 U_g826A (.Q(g826A),.SE(test_seA),.SI(g1806A),.D(g8245A),.CK(CKA));
SDFF_X1 U_g1065A (.Q(g1065A),.SE(test_seA),.SI(g826A),.D(g7242A),.CK(CKA));
SDFF_X1 U_g1887A (.Q(g1887A),.SE(test_seA),.SI(g1065A),.D(g8281A),.CK(CKA));
SDFF_X1 U_g37A (.Q(g37A),.SE(test_seA),.SI(g1887A),.D(g10724A),.CK(CKA));
SDFF_X1 U_g968A (.Q(g968A),.SE(test_seA),.SI(g37A),.D(g11314A),.CK(CKA));
SDFF_X1 U_g1845A (.Q(g1845A),.SE(test_seA),.SI(g968A),.D(g4905A),.CK(CKA));
SDFF_X1 U_g1137A (.Q(g1137A),.SE(test_seA),.SI(g1845A),.D(g4484A),.CK(CKA));
SDFF_X1 U_g1891A (.Q(g1891A),.SE(test_seA),.SI(g1137A),.D(g8937A),.CK(CKA));
SDFF_X1 U_g1255A (.Q(g1255A),.SE(test_seA),.SI(g1891A),.D(g7300A),.CK(CKA));
SDFF_X1 U_g257A (.Q(g257A),.SE(test_seA),.SI(g1255A),.D(g6002A),.CK(CKA));
SDFF_X1 U_g874A (.Q(g874A),.SE(test_seA),.SI(g257A),.D(g9507A),.CK(CKA));
SDFF_X1 U_g591A (.Q(g591A),.SE(test_seA),.SI(g874A),.D(g9110A),.CK(CKA));
SDFF_X1 U_g731A (.Q(g731A),.SE(test_seA),.SI(g591A),.D(g8926A),.CK(CKA));
SDFF_X1 U_g636A (.Q(g636A),.SE(test_seA),.SI(g731A),.D(g8631A),.CK(CKA));
SDFF_X1 U_g1218A (.Q(g1218A),.SE(test_seA),.SI(g636A),.D(g7632A),.CK(CKA));
SDFF_X1 U_g605A (.Q(g605A),.SE(test_seA),.SI(g1218A),.D(g9150A),.CK(CKA));
SDFF_X1 U_g79A (.Q(g79A),.SE(test_seA),.SI(g605A),.D(g6531A),.CK(CKA));
SDFF_X1 U_g182A (.Q(g182A),.SE(test_seA),.SI(g79A),.D(g6786A),.CK(CKA));
SDFF_X1 U_g950A (.Q(g950A),.SE(test_seA),.SI(g182A),.D(g11303A),.CK(CKA));
SDFF_X1 U_g1129A (.Q(g1129A),.SE(test_seA),.SI(g950A),.D(g4477A),.CK(CKA));
SDFF_X1 U_g857A (.Q(g857A),.SE(test_seA),.SI(g1129A),.D(g822A),.CK(CKA));
SDFF_X1 U_g448A (.Q(g448A),.SE(test_seA),.SI(g857A),.D(g11258A),.CK(CKA));
SDFF_X1 U_g1828A (.Q(g1828A),.SE(test_seA),.SI(g448A),.D(g9272A),.CK(CKA));
SDFF_X1 U_g1727A (.Q(g1727A),.SE(test_seA),.SI(g1828A),.D(g10773A),.CK(CKA));
SDFF_X1 U_g1592A (.Q(g1592A),.SE(test_seA),.SI(g1727A),.D(g6470A),.CK(CKA));
SDFF_X1 U_g1703A (.Q(g1703A),.SE(test_seA),.SI(g1592A),.D(g5083A),.CK(CKA));
SDFF_X1 U_g1932A (.Q(g1932A),.SE(test_seA),.SI(g1703A),.D(g8286A),.CK(CKA));
SDFF_X1 U_g1624A (.Q(g1624A),.SE(test_seA),.SI(g1932A),.D(g8773A),.CK(CKA));
SDFF_X1 U_g26A (.Q(g26A),.SE(test_seA),.SI(g1624A),.D(g4158A),.CK(CKA));
SDFF_X1 U_g1068A (.Q(g1068A),.SE(test_seA),.SI(g26A),.D(g6054A),.CK(CKA));
SDFF_X1 U_g578A (.Q(g578A),.SE(test_seA),.SI(g1068A),.D(g101A),.CK(CKA));
SDFF_X1 U_g440A (.Q(g440A),.SE(test_seA),.SI(g578A),.D(g11260A),.CK(CKA));
SDFF_X1 U_g476A (.Q(g476A),.SE(test_seA),.SI(g440A),.D(g11338A),.CK(CKA));
SDFF_X1 U_g119A (.Q(g119A),.SE(test_seA),.SI(g476A),.D(g5918A),.CK(CKA));
SDFF_X1 U_g668A (.Q(g668A),.SE(test_seA),.SI(g119A),.D(g8922A),.CK(CKA));
SDFF_X1 U_g139A (.Q(g139A),.SE(test_seA),.SI(g668A),.D(g8049A),.CK(CKA));
SDFF_X1 U_g1149A (.Q(g1149A),.SE(test_seA),.SI(g139A),.D(g4342A),.CK(CKA));
SDFF_X1 U_g34A (.Q(g34A),.SE(test_seA),.SI(g1149A),.D(g10720A),.CK(CKA));
SDFF_X1 U_g1848A (.Q(g1848A),.SE(test_seA),.SI(g34A),.D(g6755A),.CK(CKA));
SDFF_X1 U_g263A (.Q(g263A),.SE(test_seA),.SI(g1848A),.D(g6897A),.CK(CKA));
SDFF_X1 U_g818A (.Q(g818A),.SE(test_seA),.SI(g263A),.D(g7709A),.CK(CKA));
SDFF_X1 U_g1747A (.Q(g1747A),.SE(test_seA),.SI(g818A),.D(g4255A),.CK(CKA));
SDFF_X1 U_g802A (.Q(g802A),.SE(test_seA),.SI(g1747A),.D(g5543A),.CK(CKA));
SDFF_X1 U_g275A (.Q(g275A),.SE(test_seA),.SI(g802A),.D(g6915A),.CK(CKA));
SDFF_X1 U_g1524A (.Q(g1524A),.SE(test_seA),.SI(g275A),.D(g6513A),.CK(CKA));
SDFF_X1 U_g1577A (.Q(g1577A),.SE(test_seA),.SI(g1524A),.D(g6480A),.CK(CKA));
SDFF_X1 U_g810A (.Q(g810A),.SE(test_seA),.SI(g1577A),.D(g6733A),.CK(CKA));
SDFF_X1 U_g391A (.Q(g391A),.SE(test_seA),.SI(g810A),.D(g11264A),.CK(CKA));
SDFF_X1 U_g658A (.Q(g658A),.SE(test_seA),.SI(g391A),.D(g8973A),.CK(CKA));
SDFF_X1 U_g1386A (.Q(g1386A),.SE(test_seA),.SI(g658A),.D(g6833A),.CK(CKA));
SDFF_X1 U_g253A (.Q(g253A),.SE(test_seA),.SI(g1386A),.D(g5996A),.CK(CKA));
SDFF_X1 U_g875A (.Q(g875A),.SE(test_seA),.SI(g253A),.D(g9508A),.CK(CKA));
SDFF_X1 U_g1125A (.Q(g1125A),.SE(test_seA),.SI(g875A),.D(g4473A),.CK(CKA));
SDFF_X1 U_g201A (.Q(g201A),.SE(test_seA),.SI(g1125A),.D(g5755A),.CK(CKA));
SDFF_X1 U_g1280A (.Q(g1280A),.SE(test_seA),.SI(g201A),.D(g7295A),.CK(CKA));
SDFF_X1 U_g1083A (.Q(g1083A),.SE(test_seA),.SI(g1280A),.D(g6068A),.CK(CKA));
SDFF_X1 U_g650A (.Q(g650A),.SE(test_seA),.SI(g1083A),.D(g7137A),.CK(CKA));
SDFF_X1 U_g1636A (.Q(g1636A),.SE(test_seA),.SI(g650A),.D(g8779A),.CK(CKA));
SDFF_X1 U_g853A (.Q(g853A),.SE(test_seA),.SI(g1636A),.D(g818A),.CK(CKA));
SDFF_X1 U_g421A (.Q(g421A),.SE(test_seA),.SI(g853A),.D(g11270A),.CK(CKA));
SDFF_X1 U_g762A (.Q(g762A),.SE(test_seA),.SI(g421A),.D(g5529A),.CK(CKA));
SDFF_X1 U_g956A (.Q(g956A),.SE(test_seA),.SI(g762A),.D(g11306A),.CK(CKA));
SDFF_X1 U_g378A (.Q(g378A),.SE(test_seA),.SI(g956A),.D(g11291A),.CK(CKA));
SDFF_X1 U_g1756A (.Q(g1756A),.SE(test_seA),.SI(g378A),.D(g4283A),.CK(CKA));
SDFF_X1 U_g589A (.Q(g589A),.SE(test_seA),.SI(g1756A),.D(g29A),.CK(CKA));
SDFF_X1 U_g841A (.Q(g841A),.SE(test_seA),.SI(g589A),.D(g806A),.CK(CKA));
SDFF_X1 U_g1027A (.Q(g1027A),.SE(test_seA),.SI(g841A),.D(g6894A),.CK(CKA));
SDFF_X1 U_g1003A (.Q(g1003A),.SE(test_seA),.SI(g1027A),.D(g6902A),.CK(CKA));
SDFF_X1 U_g1403A (.Q(g1403A),.SE(test_seA),.SI(g1003A),.D(g8765A),.CK(CKA));
SDFF_X1 U_g1145A (.Q(g1145A),.SE(test_seA),.SI(g1403A),.D(g4498A),.CK(CKA));
SDFF_X1 U_g1107A (.Q(g1107A),.SE(test_seA),.SI(g1145A),.D(g5148A),.CK(CKA));
SDFF_X1 U_g1223A (.Q(g1223A),.SE(test_seA),.SI(g1107A),.D(g7581A),.CK(CKA));
SDFF_X1 U_g406A (.Q(g406A),.SE(test_seA),.SI(g1223A),.D(g11267A),.CK(CKA));
SDFF_X1 U_g1811A (.Q(g1811A),.SE(test_seA),.SI(g406A),.D(g10936A),.CK(CKA));
SDFF_X1 U_g1642A (.Q(g1642A),.SE(test_seA),.SI(g1811A),.D(g10784A),.CK(CKA));
SDFF_X1 U_g1047A (.Q(g1047A),.SE(test_seA),.SI(g1642A),.D(g7211A),.CK(CKA));
SDFF_X1 U_g1654A (.Q(g1654A),.SE(test_seA),.SI(g1047A),.D(g10765A),.CK(CKA));
SDFF_X1 U_g197A (.Q(g197A),.SE(test_seA),.SI(g1654A),.D(g6332A),.CK(CKA));
SDFF_X1 U_g1595A (.Q(g1595A),.SE(test_seA),.SI(g197A),.D(g6479A),.CK(CKA));
SDFF_X1 U_g1537A (.Q(g1537A),.SE(test_seA),.SI(g1595A),.D(g6537A),.CK(CKA));
SDFF_X1 U_g727A (.Q(g727A),.SE(test_seA),.SI(g1537A),.D(g8434A),.CK(CKA));
SDFF_X1 U_g999A (.Q(g999A),.SE(test_seA),.SI(g727A),.D(g6908A),.CK(CKA));
SDFF_X1 U_g798A (.Q(g798A),.SE(test_seA),.SI(g999A),.D(g6243A),.CK(CKA));
SDFF_X1 U_g481A (.Q(g481A),.SE(test_seA),.SI(g798A),.D(g11324A),.CK(CKA));
SDFF_X1 U_g754A (.Q(g754A),.SE(test_seA),.SI(g481A),.D(g3462A),.CK(CKA));
SDFF_X1 U_g1330A (.Q(g1330A),.SE(test_seA),.SI(g754A),.D(g11609A),.CK(CKA));
SDFF_X1 U_g845A (.Q(g845A),.SE(test_seA),.SI(g1330A),.D(g810A),.CK(CKA));
SDFF_X1 U_g790A (.Q(g790A),.SE(test_seA),.SI(g845A),.D(g8244A),.CK(CKA));
SDFF_X1 U_g1512A (.Q(g1512A),.SE(test_seA),.SI(g790A),.D(g8194A),.CK(CKA));
SDFF_X1 U_g114A (.Q(g114A),.SE(test_seA),.SI(g1512A),.D(g113A),.CK(CKA));
SDFF_X1 U_g1490A (.Q(g1490A),.SE(test_seA),.SI(g114A),.D(g8052A),.CK(CKA));
SDFF_X1 U_g1166A (.Q(g1166A),.SE(test_seA),.SI(g1490A),.D(g4325A),.CK(CKA));
SDFF_X1 U_g1056A (.Q(g1056A),.SE(test_seA),.SI(g1166A),.D(g7231A),.CK(CKA));
SDFF_X1 U_g348A (.Q(g348A),.SE(test_seA),.SI(g1056A),.D(g11481A),.CK(CKA));
SDFF_X1 U_g868A (.Q(g868A),.SE(test_seA),.SI(g348A),.D(g874A),.CK(CKA));
SDFF_X1 U_g1260A (.Q(g1260A),.SE(test_seA),.SI(g868A),.D(g7301A),.CK(CKA));
SDFF_X1 U_g260A (.Q(g260A),.SE(test_seA),.SI(g1260A),.D(g6035A),.CK(CKA));
SDFF_X1 U_g131A (.Q(g131A),.SE(test_seA),.SI(g260A),.D(g8059A),.CK(CKA));
SDFF_X1 U_g7A (.Q(g7A),.SE(test_seA),.SI(g131A),.D(g1854A),.CK(CKA));
SDFF_X1 U_g258A (.Q(g258A),.SE(test_seA),.SI(g7A),.D(g6015A),.CK(CKA));
SDFF_X1 U_g521A (.Q(g521A),.SE(test_seA),.SI(g258A),.D(g11330A),.CK(CKA));
SDFF_X1 U_g1318A (.Q(g1318A),.SE(test_seA),.SI(g521A),.D(g11605A),.CK(CKA));
SDFF_X1 U_g1872A (.Q(g1872A),.SE(test_seA),.SI(g1318A),.D(g8921A),.CK(CKA));
SDFF_X1 U_g677A (.Q(g677A),.SE(test_seA),.SI(g1872A),.D(g8883A),.CK(CKA));
SDFF_X1 U_g582A (.Q(g582A),.SE(test_seA),.SI(g677A),.D(g28A),.CK(CKA));
SDFF_X1 U_g1393A (.Q(g1393A),.SE(test_seA),.SI(g582A),.D(g6163A),.CK(CKA));
SDFF_X1 U_g1549A (.Q(g1549A),.SE(test_seA),.SI(g1393A),.D(g6523A),.CK(CKA));
SDFF_X1 U_g947A (.Q(g947A),.SE(test_seA),.SI(g1549A),.D(g11300A),.CK(CKA));
SDFF_X1 U_g1834A (.Q(g1834A),.SE(test_seA),.SI(g947A),.D(g9555A),.CK(CKA));
SDFF_X1 U_g1598A (.Q(g1598A),.SE(test_seA),.SI(g1834A),.D(g6481A),.CK(CKA));
SDFF_X1 U_g1121A (.Q(g1121A),.SE(test_seA),.SI(g1598A),.D(g4471A),.CK(CKA));
SDFF_X1 U_g1321A (.Q(g1321A),.SE(test_seA),.SI(g1121A),.D(g11606A),.CK(CKA));
SDFF_X1 U_g506A (.Q(g506A),.SE(test_seA),.SI(g1321A),.D(g11335A),.CK(CKA));
SDFF_X1 U_g546A (.Q(g546A),.SE(test_seA),.SI(g506A),.D(g10791A),.CK(CKA));
SDFF_X1 U_g1909A (.Q(g1909A),.SE(test_seA),.SI(g546A),.D(g8939A),.CK(CKA));
SDFF_X1 U_g755A (.Q(g755A),.SE(test_seA),.SI(g1909A),.D(g83A),.CK(CKA));
SDFF_X1 U_g1552A (.Q(g1552A),.SE(test_seA),.SI(g755A),.D(g6529A),.CK(CKA));
SDFF_X1 U_g584A (.Q(g584A),.SE(test_seA),.SI(g1552A),.D(g101A),.CK(CKA));
SDFF_X1 U_g1687A (.Q(g1687A),.SE(test_seA),.SI(g584A),.D(g10776A),.CK(CKA));
SDFF_X1 U_g1586A (.Q(g1586A),.SE(test_seA),.SI(g1687A),.D(g6514A),.CK(CKA));
SDFF_X1 U_g324A (.Q(g324A),.SE(test_seA),.SI(g1586A),.D(g259A),.CK(CKA));
SDFF_X1 U_g1141A (.Q(g1141A),.SE(test_seA),.SI(g324A),.D(g4490A),.CK(CKA));
SDFF_X1 U_g1570A (.Q(g1570A),.SE(test_seA),.SI(g1141A),.D(I8503A),.CK(CKA));
SDFF_X1 U_g1341A (.Q(g1341A),.SE(test_seA),.SI(g1570A),.D(g11639A),.CK(CKA));
SDFF_X1 U_g1710A (.Q(g1710A),.SE(test_seA),.SI(g1341A),.D(g4089A),.CK(CKA));
SDFF_X1 U_g1645A (.Q(g1645A),.SE(test_seA),.SI(g1710A),.D(g10785A),.CK(CKA));
SDFF_X1 U_g115A (.Q(g115A),.SE(test_seA),.SI(g1645A),.D(g6179A),.CK(CKA));
SDFF_X1 U_g135A (.Q(g135A),.SE(test_seA),.SI(g115A),.D(g8053A),.CK(CKA));
SDFF_X1 U_g525A (.Q(g525A),.SE(test_seA),.SI(g135A),.D(g11329A),.CK(CKA));
SDFF_X1 U_g581A (.Q(g581A),.SE(test_seA),.SI(g525A),.D(g104A),.CK(CKA));
SDFF_X1 U_g1607A (.Q(g1607A),.SE(test_seA),.SI(g581A),.D(g6515A),.CK(CKA));
SDFF_X1 U_g321A (.Q(g321A),.SE(test_seA),.SI(g1607A),.D(g258A),.CK(CKA));
SDFF_X1 U_g67A (.Q(g67A),.SE(test_seA),.SI(g321A),.D(g7204A),.CK(CKA));
SDFF_X1 U_g1275A (.Q(g1275A),.SE(test_seA),.SI(g67A),.D(g11443A),.CK(CKA));
SDFF_X1 U_g1311A (.Q(g1311A),.SE(test_seA),.SI(g1275A),.D(g11603A),.CK(CKA));
SDFF_X1 U_g1615A (.Q(g1615A),.SE(test_seA),.SI(g1311A),.D(g8770A),.CK(CKA));
SDFF_X1 U_g382A (.Q(g382A),.SE(test_seA),.SI(g1615A),.D(g11292A),.CK(CKA));
SDFF_X1 U_g1374A (.Q(g1374A),.SE(test_seA),.SI(g382A),.D(g6331A),.CK(CKA));
SDFF_X1 U_g266A (.Q(g266A),.SE(test_seA),.SI(g1374A),.D(g6900A),.CK(CKA));
SDFF_X1 U_g1284A (.Q(g1284A),.SE(test_seA),.SI(g266A),.D(g7294A),.CK(CKA));
SDFF_X1 U_g1380A (.Q(g1380A),.SE(test_seA),.SI(g1284A),.D(g6829A),.CK(CKA));
SDFF_X1 U_g673A (.Q(g673A),.SE(test_seA),.SI(g1380A),.D(g8428A),.CK(CKA));
SDFF_X1 U_g1853A (.Q(g1853A),.SE(test_seA),.SI(g673A),.D(g4904A),.CK(CKA));
SDFF_X1 U_g162A (.Q(g162A),.SE(test_seA),.SI(g1853A),.D(g8054A),.CK(CKA));
SDFF_X1 U_g411A (.Q(g411A),.SE(test_seA),.SI(g162A),.D(g11268A),.CK(CKA));
SDFF_X1 U_g431A (.Q(g431A),.SE(test_seA),.SI(g411A),.D(g11262A),.CK(CKA));
SDFF_X1 U_g1905A (.Q(g1905A),.SE(test_seA),.SI(g431A),.D(g8283A),.CK(CKA));
SDFF_X1 U_g1515A (.Q(g1515A),.SE(test_seA),.SI(g1905A),.D(g6193A),.CK(CKA));
SDFF_X1 U_g1630A (.Q(g1630A),.SE(test_seA),.SI(g1515A),.D(g8776A),.CK(CKA));
SDFF_X1 U_g49A (.Q(g49A),.SE(test_seA),.SI(g1630A),.D(g7143A),.CK(CKA));
SDFF_X1 U_g991A (.Q(g991A),.SE(test_seA),.SI(g49A),.D(g6898A),.CK(CKA));
SDFF_X1 U_g1300A (.Q(g1300A),.SE(test_seA),.SI(g991A),.D(g7291A),.CK(CKA));
SDFF_X1 U_g339A (.Q(g339A),.SE(test_seA),.SI(g1300A),.D(g11478A),.CK(CKA));
SDFF_X1 U_g256A (.Q(g256A),.SE(test_seA),.SI(g339A),.D(g6000A),.CK(CKA));
SDFF_X1 U_g1750A (.Q(g1750A),.SE(test_seA),.SI(g256A),.D(g4264A),.CK(CKA));
SDFF_X1 U_g585A (.Q(g585A),.SE(test_seA),.SI(g1750A),.D(g102A),.CK(CKA));
SDFF_X1 U_g1440A (.Q(g1440A),.SE(test_seA),.SI(g585A),.D(g8768A),.CK(CKA));
SDFF_X1 U_g1666A (.Q(g1666A),.SE(test_seA),.SI(g1440A),.D(g10863A),.CK(CKA));
SDFF_X1 U_g1528A (.Q(g1528A),.SE(test_seA),.SI(g1666A),.D(g6522A),.CK(CKA));
SDFF_X1 U_g1351A (.Q(g1351A),.SE(test_seA),.SI(g1528A),.D(g11641A),.CK(CKA));
SDFF_X1 U_g1648A (.Q(g1648A),.SE(test_seA),.SI(g1351A),.D(g10780A),.CK(CKA));
SDFF_X1 U_g127A (.Q(g127A),.SE(test_seA),.SI(g1648A),.D(g8044A),.CK(CKA));
SDFF_X1 U_g1618A (.Q(g1618A),.SE(test_seA),.SI(g127A),.D(g11579A),.CK(CKA));
SDFF_X1 U_g1235A (.Q(g1235A),.SE(test_seA),.SI(g1618A),.D(g7296A),.CK(CKA));
SDFF_X1 U_g299A (.Q(g299A),.SE(test_seA),.SI(g1235A),.D(g6923A),.CK(CKA));
SDFF_X1 U_g435A (.Q(g435A),.SE(test_seA),.SI(g299A),.D(g11261A),.CK(CKA));
SDFF_X1 U_g64A (.Q(g64A),.SE(test_seA),.SI(g435A),.D(g6638A),.CK(CKA));
SDFF_X1 U_g1555A (.Q(g1555A),.SE(test_seA),.SI(g64A),.D(g6534A),.CK(CKA));
SDFF_X1 U_g995A (.Q(g995A),.SE(test_seA),.SI(g1555A),.D(g6895A),.CK(CKA));
SDFF_X1 U_g1621A (.Q(g1621A),.SE(test_seA),.SI(g995A),.D(g8771A),.CK(CKA));
SDFF_X1 U_g1113A (.Q(g1113A),.SE(test_seA),.SI(g1621A),.D(g4506A),.CK(CKA));
SDFF_X1 U_g643A (.Q(g643A),.SE(test_seA),.SI(g1113A),.D(g7441A),.CK(CKA));
SDFF_X1 U_g1494A (.Q(g1494A),.SE(test_seA),.SI(g643A),.D(g8055A),.CK(CKA));
SDFF_X1 U_g1567A (.Q(g1567A),.SE(test_seA),.SI(g1494A),.D(g6468A),.CK(CKA));
SDFF_X1 U_g691A (.Q(g691A),.SE(test_seA),.SI(g1567A),.D(g8430A),.CK(CKA));
SDFF_X1 U_g534A (.Q(g534A),.SE(test_seA),.SI(g691A),.D(g11327A),.CK(CKA));
SDFF_X1 U_g1776A (.Q(g1776A),.SE(test_seA),.SI(g534A),.D(g6508A),.CK(CKA));
SDFF_X1 U_g569A (.Q(g569A),.SE(test_seA),.SI(g1776A),.D(g10717A),.CK(CKA));
SDFF_X1 U_g1160A (.Q(g1160A),.SE(test_seA),.SI(g569A),.D(g4334A),.CK(CKA));
SDFF_X1 U_g1360A (.Q(g1360A),.SE(test_seA),.SI(g1160A),.D(g9526A),.CK(CKA));
SDFF_X1 U_g1050A (.Q(g1050A),.SE(test_seA),.SI(g1360A),.D(g7218A),.CK(CKA));
SDFF_X1 U_g1A (.Q(g1A),.SE(test_seA),.SI(g1050A),.D(g6679A),.CK(CKA));
SDFF_X1 U_g511A (.Q(g511A),.SE(test_seA),.SI(g1A),.D(g11336A),.CK(CKA));
SDFF_X1 U_g1724A (.Q(g1724A),.SE(test_seA),.SI(g511A),.D(g10771A),.CK(CKA));
SDFF_X1 U_g12A (.Q(g12A),.SE(test_seA),.SI(g1724A),.D(g5445A),.CK(CKA));
SDFF_X1 U_g1878A (.Q(g1878A),.SE(test_seA),.SI(g12A),.D(g8559A),.CK(CKA));
SDFF_X1 U_g73A (.Q(g73A),.SE(test_seA),.SI(g1878A),.D(g7219A),.CK(CKA));
INV_X1 FE_OFC370_g4525B (.ZN(FE_OFN370_g4525B),.A(FE_OFN368_g4525B));
INV_X1 FE_OFC369_g4525B (.ZN(FE_OFN369_g4525B),.A(FE_OFN368_g4525B));
INV_X1 FE_OFC368_g4525B (.ZN(FE_OFN368_g4525B),.A(FE_OFN362_g4525B));
BUF_X3 FE_OFC367_g3521B (.Z(FE_OFN367_g3521B),.A(FE_OFN366_g3521B));
BUF_X3 FE_OFC366_g3521B (.Z(FE_OFN366_g3521B),.A(FE_OFN358_g3521B));
BUF_X3 FE_OFC365_g5361B (.Z(FE_OFN365_g5361B),.A(FE_OFN356_g5361B));
BUF_X3 FE_OFC364_g3015B (.Z(FE_OFN364_g3015B),.A(FE_OFN348_g3015B));
BUF_X3 FE_OFC363_I5565B (.Z(FE_OFN363_I5565B),.A(FE_OFN343_I5565B));
INV_X1 FE_OFC362_g4525B (.ZN(FE_OFN362_g4525B),.A(FE_OFN360_g4525B));
INV_X1 FE_OFC360_g4525B (.ZN(FE_OFN360_g4525B),.A(FE_OFN339_g4525B));
BUF_X3 FE_OFC359_g18B (.Z(FE_OFN359_g18B),.A(FE_OFN324_g18B));
BUF_X3 FE_OFC358_g3521B (.Z(FE_OFN358_g3521B),.A(g3521B));
BUF_X3 FE_OFC357_g3521B (.Z(FE_OFN357_g3521B),.A(FE_OFN366_g3521B));
INV_X1 FE_OFC356_g5361B (.ZN(FE_OFN356_g5361B),.A(FE_OFN354_g5361B));
INV_X1 FE_OFC354_g5361B (.ZN(FE_OFN354_g5361B),.A(FE_OFN318_g5361B));
BUF_X3 FE_OFC353_g5117B (.Z(FE_OFN353_g5117B),.A(FE_OFN315_g5117B));
BUF_X3 FE_OFC352_g109B (.Z(FE_OFN352_g109B),.A(FE_OFN269_g109B));
BUF_X3 FE_OFC351_g3913B (.Z(FE_OFN351_g3913B),.A(FE_OFN302_g3913B));
BUF_X3 FE_OFC350_g3121B (.Z(FE_OFN350_g3121B),.A(FE_OFN155_g3121B));
BUF_X3 FE_OFC349_I6424B (.Z(FE_OFN349_I6424B),.A(FE_OFN308_I6424B));
BUF_X3 FE_OFC348_g3015B (.Z(FE_OFN348_g3015B),.A(FE_OFN298_g3015B));
BUF_X3 FE_OFC347_g3914B (.Z(FE_OFN347_g3914B),.A(FE_OFN296_g3914B));
BUF_X3 FE_OFC346_g4381B (.Z(FE_OFN346_g4381B),.A(g4381B));
BUF_X3 FE_OFC345_g3015B (.Z(FE_OFN345_g3015B),.A(FE_OFN297_g3015B));
BUF_X3 FE_OFC344_g3586B (.Z(FE_OFN344_g3586B),.A(FE_OFN287_g3586B));
INV_X1 FE_OFC343_I5565B (.ZN(FE_OFN343_I5565B),.A(FE_OFN340_I5565B));
INV_X1 FE_OFC340_I5565B (.ZN(FE_OFN340_I5565B),.A(FE_OFN233_I5565B));
INV_X1 FE_OFC339_g4525B (.ZN(FE_OFN339_g4525B),.A(FE_OFN337_g4525B));
INV_X1 FE_OFC337_g4525B (.ZN(FE_OFN337_g4525B),.A(g4525B));
BUF_X3 FE_OFC336_g1690B (.Z(FE_OFN336_g1690B),.A(FE_OFN245_g1690B));
BUF_X3 FE_OFC335_g4737B (.Z(FE_OFN335_g4737B),.A(g4737B));
BUF_X3 FE_OFC334_g7045B (.Z(FE_OFN334_g7045B),.A(g7045B));
BUF_X3 FE_OFC333_g4294B (.Z(FE_OFN333_g4294B),.A(g4294B));
BUF_X3 FE_OFC332_g8748B (.Z(FE_OFN332_g8748B),.A(g8748B));
BUF_X3 FE_OFC331_g8696B (.Z(FE_OFN331_g8696B),.A(g8696B));
BUF_X3 FE_OFC330_g7638B (.Z(FE_OFN330_g7638B),.A(FE_OFN189_g7638B));
BUF_X3 FE_OFC329_g8763B (.Z(FE_OFN329_g8763B),.A(g8763B));
BUF_X3 FE_OFC328_g8709B (.Z(FE_OFN328_g8709B),.A(g8709B));
BUF_X3 FE_OFC325_g18B (.Z(FE_OFN325_g18B),.A(FE_OFN359_g18B));
BUF_X3 FE_OFC324_g18B (.Z(FE_OFN324_g18B),.A(FE_OFN260_g18B));
BUF_X3 FE_OFC322_g4449B (.Z(FE_OFN322_g4449B),.A(g4449B));
BUF_X3 FE_OFC321_g5261B (.Z(FE_OFN321_g5261B),.A(g5261B));
BUF_X3 FE_OFC320_g5361B (.Z(FE_OFN320_g5361B),.A(FE_OFN319_g5361B));
BUF_X3 FE_OFC319_g5361B (.Z(FE_OFN319_g5361B),.A(FE_OFN166_g5361B));
INV_X1 FE_OFC318_g5361B (.ZN(FE_OFN318_g5361B),.A(FE_OFN316_g5361B));
INV_X1 FE_OFC316_g5361B (.ZN(FE_OFN316_g5361B),.A(FE_OFN168_g5361B));
INV_X1 FE_OFC315_g5117B (.ZN(FE_OFN315_g5117B),.A(FE_OFN312_g5117B));
INV_X1 FE_OFC312_g5117B (.ZN(FE_OFN312_g5117B),.A(g5117B));
BUF_X3 FE_OFC310_g4336B (.Z(FE_OFN310_g4336B),.A(g4336B));
BUF_X3 FE_OFC308_I6424B (.Z(FE_OFN308_I6424B),.A(FE_OFN160_I6424B));
BUF_X3 FE_OFC307_g4010B (.Z(FE_OFN307_g4010B),.A(g4010B));
BUF_X3 FE_OFC306_g5128B (.Z(FE_OFN306_g5128B),.A(g5128B));
BUF_X3 FE_OFC305_g5151B (.Z(FE_OFN305_g5151B),.A(FE_OFN304_g5151B));
BUF_X3 FE_OFC304_g5151B (.Z(FE_OFN304_g5151B),.A(FE_OFN176_g5151B));
BUF_X3 FE_OFC303_g4678B (.Z(FE_OFN303_g4678B),.A(g4678B));
BUF_X3 FE_OFC302_g3913B (.Z(FE_OFN302_g3913B),.A(g3913B));
BUF_X3 FE_OFC300_g4002B (.Z(FE_OFN300_g4002B),.A(g4002B));
BUF_X3 FE_OFC299_g4457B (.Z(FE_OFN299_g4457B),.A(g4457B));
BUF_X3 FE_OFC298_g3015B (.Z(FE_OFN298_g3015B),.A(FE_OFN119_g3015B));
BUF_X3 FE_OFC297_g3015B (.Z(FE_OFN297_g3015B),.A(FE_OFN348_g3015B));
INV_X1 FE_OFC296_g3914B (.ZN(FE_OFN296_g3914B),.A(FE_OFN294_g3914B));
INV_X1 FE_OFC294_g3914B (.ZN(FE_OFN294_g3914B),.A(FE_OFN113_g3914B));
BUF_X3 FE_OFC293_g3015B (.Z(FE_OFN293_g3015B),.A(FE_OFN292_g3015B));
BUF_X3 FE_OFC292_g3015B (.Z(FE_OFN292_g3015B),.A(FE_OFN345_g3015B));
BUF_X3 FE_OFC291_g4880B (.Z(FE_OFN291_g4880B),.A(FE_OFN290_g4880B));
BUF_X3 FE_OFC290_g4880B (.Z(FE_OFN290_g4880B),.A(g4880B));
BUF_X3 FE_OFC289_g4679B (.Z(FE_OFN289_g4679B),.A(g4679B));
BUF_X3 FE_OFC288_g4263B (.Z(FE_OFN288_g4263B),.A(g4263B));
INV_X1 FE_OFC287_g3586B (.ZN(FE_OFN287_g3586B),.A(FE_OFN284_g3586B));
INV_X1 FE_OFC284_g3586B (.ZN(FE_OFN284_g3586B),.A(FE_OFN110_g3586B));
BUF_X3 FE_OFC283_I8869B (.Z(FE_OFN283_I8869B),.A(FE_OFN97_I8869B));
BUF_X3 FE_OFC282_g6165B (.Z(FE_OFN282_g6165B),.A(g6165B));
BUF_X3 FE_OFC281_g2216B (.Z(FE_OFN281_g2216B),.A(FE_OFN95_g2216B));
BUF_X3 FE_OFC280_g9536B (.Z(FE_OFN280_g9536B),.A(FE_OFN64_g9536B));
BUF_X3 FE_OFC279_g11157B (.Z(FE_OFN279_g11157B),.A(g11157B));
BUF_X3 FE_OFC278_g10927B (.Z(FE_OFN278_g10927B),.A(g10927B));
BUF_X3 FE_OFC277_g48B (.Z(FE_OFN277_g48B),.A(FE_OFN276_g48B));
BUF_X3 FE_OFC276_g48B (.Z(FE_OFN276_g48B),.A(FE_OFN275_g48B));
BUF_X3 FE_OFC275_g48B (.Z(FE_OFN275_g48B),.A(g48B));
BUF_X3 FE_OFC273_g85B (.Z(FE_OFN273_g85B),.A(FE_OFN271_g85B));
BUF_X3 FE_OFC271_g85B (.Z(FE_OFN271_g85B),.A(g85B));
BUF_X3 FE_OFC269_g109B (.Z(FE_OFN269_g109B),.A(FE_OFN267_g109B));
BUF_X3 FE_OFC267_g109B (.Z(FE_OFN267_g109B),.A(g109B));
BUF_X3 FE_OFC266_g18B (.Z(FE_OFN266_g18B),.A(FE_OFN325_g18B));
BUF_X3 FE_OFC260_g18B (.Z(FE_OFN260_g18B),.A(g2355B));
BUF_X3 FE_OFC254_g461B (.Z(FE_OFN254_g461B),.A(g461B));
BUF_X3 FE_OFC253_g1786B (.Z(FE_OFN253_g1786B),.A(g1786B));
BUF_X3 FE_OFC252_g1791B (.Z(FE_OFN252_g1791B),.A(g1791B));
BUF_X3 FE_OFC251_g1801B (.Z(FE_OFN251_g1801B),.A(g1801B));
BUF_X3 FE_OFC250_g471B (.Z(FE_OFN250_g471B),.A(g471B));
BUF_X3 FE_OFC248_g466B (.Z(FE_OFN248_g466B),.A(g466B));
BUF_X3 FE_OFC247_g1771B (.Z(FE_OFN247_g1771B),.A(g1771B));
INV_X1 FE_OFC245_g1690B (.ZN(FE_OFN245_g1690B),.A(g2424B));
BUF_X3 FE_OFC241_g1690B (.Z(FE_OFN241_g1690B),.A(g1690B));
BUF_X3 FE_OFC240_g1110B (.Z(FE_OFN240_g1110B),.A(g1110B));
BUF_X3 FE_OFC239_g1796B (.Z(FE_OFN239_g1796B),.A(g1796B));
BUF_X3 FE_OFC238_g1781B (.Z(FE_OFN238_g1781B),.A(g1781B));
BUF_X3 FE_OFC237_g1806B (.Z(FE_OFN237_g1806B),.A(g1806B));
BUF_X3 FE_OFC236_g1776B (.Z(FE_OFN236_g1776B),.A(g1776B));
BUF_X3 FE_OFC235_g2024B (.Z(FE_OFN235_g2024B),.A(FE_OFN234_g2024B));
BUF_X3 FE_OFC234_g2024B (.Z(FE_OFN234_g2024B),.A(g2024B));
INV_X1 FE_OFC233_I5565B (.ZN(FE_OFN233_I5565B),.A(FE_OFN230_I5565B));
INV_X1 FE_OFC230_I5565B (.ZN(FE_OFN230_I5565B),.A(I6360B));
INV_X1 FE_OFC229_g3880B (.ZN(FE_OFN229_g3880B),.A(FE_OFN227_g3880B));
INV_X1 FE_OFC227_g3880B (.ZN(FE_OFN227_g3880B),.A(FE_OFN226_g3880B));
BUF_X3 FE_OFC226_g3880B (.Z(FE_OFN226_g3880B),.A(g3880B));
BUF_X3 FE_OFC225_g2276B (.Z(FE_OFN225_g2276B),.A(FE_OFN224_g2276B));
BUF_X3 FE_OFC224_g2276B (.Z(FE_OFN224_g2276B),.A(g2276B));
BUF_X3 FE_OFC223_g4401B (.Z(FE_OFN223_g4401B),.A(g4401B));
BUF_X3 FE_OFC221_g3440B (.Z(FE_OFN221_g3440B),.A(g3440B));
BUF_X3 FE_OFC219_g5557B (.Z(FE_OFN219_g5557B),.A(FE_OFN218_g5557B));
BUF_X3 FE_OFC218_g5557B (.Z(FE_OFN218_g5557B),.A(g5557B));
INV_X1 FE_OFC217_g5013B (.ZN(FE_OFN217_g5013B),.A(g6403B));
BUF_X3 FE_OFC213_g6003B (.Z(FE_OFN213_g6003B),.A(g6003B));
BUF_X3 FE_OFC211_g7246B (.Z(FE_OFN211_g7246B),.A(FE_OFN210_g7246B));
BUF_X3 FE_OFC210_g7246B (.Z(FE_OFN210_g7246B),.A(g7246B));
INV_X1 FE_OFC209_g6863B (.ZN(FE_OFN209_g6863B),.A(FE_OFN207_g6863B));
INV_X1 FE_OFC207_g6863B (.ZN(FE_OFN207_g6863B),.A(FE_OFN206_g6863B));
BUF_X3 FE_OFC206_g6863B (.Z(FE_OFN206_g6863B),.A(g6863B));
BUF_X3 FE_OFC204_g3664B (.Z(FE_OFN204_g3664B),.A(g3664B));
BUF_X3 FE_OFC200_g4921B (.Z(FE_OFN200_g4921B),.A(g4921B));
BUF_X3 FE_OFC199_g7697B (.Z(FE_OFN199_g7697B),.A(FE_OFN198_g7697B));
INV_X1 FE_OFC198_g7697B (.ZN(FE_OFN198_g7697B),.A(FE_OFN196_g7697B));
INV_X1 FE_OFC196_g7697B (.ZN(FE_OFN196_g7697B),.A(g7697B));
INV_X1 FE_OFC195_g6488B (.ZN(FE_OFN195_g6488B),.A(FE_OFN192_g6488B));
INV_X1 FE_OFC192_g6488B (.ZN(FE_OFN192_g6488B),.A(g6488B));
BUF_X3 FE_OFC191_g6488B (.Z(FE_OFN191_g6488B),.A(g6488B));
INV_X1 FE_OFC189_g7638B (.ZN(FE_OFN189_g7638B),.A(FE_OFN187_g7638B));
INV_X1 FE_OFC187_g7638B (.ZN(FE_OFN187_g7638B),.A(g7638B));
BUF_X3 FE_OFC184_I7048B (.Z(FE_OFN184_I7048B),.A(I7048B));
BUF_X3 FE_OFC180_g5354B (.Z(FE_OFN180_g5354B),.A(FE_OFN179_g5354B));
BUF_X3 FE_OFC179_g5354B (.Z(FE_OFN179_g5354B),.A(FE_OFN178_g5354B));
BUF_X3 FE_OFC178_g5354B (.Z(FE_OFN178_g5354B),.A(g5354B));
BUF_X3 FE_OFC177_g5919B (.Z(FE_OFN177_g5919B),.A(g5919B));
BUF_X3 FE_OFC176_g5151B (.Z(FE_OFN176_g5151B),.A(FE_OFN306_g5128B));
INV_X1 FE_OFC168_g5361B (.ZN(FE_OFN168_g5361B),.A(FE_OFN166_g5361B));
INV_X1 FE_OFC166_g5361B (.ZN(FE_OFN166_g5361B),.A(FE_OFN164_g5361B));
INV_X1 FE_OFC164_g5361B (.ZN(FE_OFN164_g5361B),.A(FE_OFN161_g5361B));
INV_X1 FE_OFC161_g5361B (.ZN(FE_OFN161_g5361B),.A(g5361B));
BUF_X3 FE_OFC160_I6424B (.Z(FE_OFN160_I6424B),.A(FE_OFN350_g3121B));
BUF_X3 FE_OFC155_g3121B (.Z(FE_OFN155_g3121B),.A(g3121B));
BUF_X3 FE_OFC154_g4640B (.Z(FE_OFN154_g4640B),.A(FE_OFN153_g4640B));
INV_X1 FE_OFC153_g4640B (.ZN(FE_OFN153_g4640B),.A(FE_OFN321_g5261B));
BUF_X4 FE_OFC147_g4682B (.Z(FE_OFN147_g4682B),.A(FE_OFN146_g4682B));
BUF_X3 FE_OFC146_g4682B (.Z(FE_OFN146_g4682B),.A(FE_OFN144_g4682B));
INV_X1 FE_OFC144_g4682B (.ZN(FE_OFN144_g4682B),.A(FE_OFN142_g4682B));
INV_X1 FE_OFC142_g4682B (.ZN(FE_OFN142_g4682B),.A(g4682B));
INV_X1 FE_OFC141_g3829B (.ZN(FE_OFN141_g3829B),.A(FE_OFN299_g4457B));
BUF_X3 FE_OFC137_g3829B (.Z(FE_OFN137_g3829B),.A(g3829B));
INV_X1 FE_OFC136_g3863B (.ZN(FE_OFN136_g3863B),.A(FE_OFN134_g3863B));
INV_X1 FE_OFC134_g3863B (.ZN(FE_OFN134_g3863B),.A(g3863B));
BUF_X3 FE_OFC133_g3015B (.Z(FE_OFN133_g3015B),.A(FE_OFN131_g3015B));
BUF_X3 FE_OFC132_g3015B (.Z(FE_OFN132_g3015B),.A(FE_OFN293_g3015B));
INV_X1 FE_OFC131_g3015B (.ZN(FE_OFN131_g3015B),.A(FE_OFN291_g4880B));
BUF_X3 FE_OFC119_g3015B (.Z(FE_OFN119_g3015B),.A(g3015B));
BUF_X3 FE_OFC118_g4807B (.Z(FE_OFN118_g4807B),.A(FE_OFN117_g4807B));
BUF_X3 FE_OFC117_g4807B (.Z(FE_OFN117_g4807B),.A(FE_OFN116_g4807B));
BUF_X3 FE_OFC116_g4807B (.Z(FE_OFN116_g4807B),.A(FE_OFN115_g4807B));
BUF_X3 FE_OFC115_g4807B (.Z(FE_OFN115_g4807B),.A(g4807B));
INV_X1 FE_OFC113_g3914B (.ZN(FE_OFN113_g3914B),.A(FE_OFN111_g3914B));
INV_X1 FE_OFC111_g3914B (.ZN(FE_OFN111_g3914B),.A(g4673B));
INV_X1 FE_OFC110_g3586B (.ZN(FE_OFN110_g3586B),.A(g4263B));
BUF_X3 FE_OFC103_g3586B (.Z(FE_OFN103_g3586B),.A(FE_OFN102_g3586B));
BUF_X3 FE_OFC102_g3586B (.Z(FE_OFN102_g3586B),.A(g3586B));
BUF_X3 FE_OFC100_g4421B (.Z(FE_OFN100_g4421B),.A(FE_OFN99_g4421B));
BUF_X3 FE_OFC99_g4421B (.Z(FE_OFN99_g4421B),.A(g4421B));
BUF_X3 FE_OFC97_I8869B (.Z(FE_OFN97_I8869B),.A(I8869B));
BUF_X3 FE_OFC96_g2169B (.Z(FE_OFN96_g2169B),.A(g2169B));
BUF_X3 FE_OFC95_g2216B (.Z(FE_OFN95_g2216B),.A(FE_OFN93_g2216B));
BUF_X3 FE_OFC93_g2216B (.Z(FE_OFN93_g2216B),.A(FE_OFN92_g2216B));
BUF_X3 FE_OFC92_g2216B (.Z(FE_OFN92_g2216B),.A(g2216B));
BUF_X3 FE_OFC91_g2172B (.Z(FE_OFN91_g2172B),.A(g2172B));
BUF_X3 FE_OFC90_I11360B (.Z(FE_OFN90_I11360B),.A(FE_OFN89_I11360B));
BUF_X3 FE_OFC89_I11360B (.Z(FE_OFN89_I11360B),.A(I11360B));
BUF_X3 FE_OFC88_g2178B (.Z(FE_OFN88_g2178B),.A(g2178B));
BUF_X3 FE_OFC87_g2176B (.Z(FE_OFN87_g2176B),.A(FE_OFN86_g2176B));
BUF_X3 FE_OFC86_g2176B (.Z(FE_OFN86_g2176B),.A(FE_OFN85_g2176B));
BUF_X3 FE_OFC85_g2176B (.Z(FE_OFN85_g2176B),.A(FE_OFN83_g2176B));
INV_X1 FE_OFC84_g2176B (.ZN(FE_OFN84_g2176B),.A(FE_OFN81_g2176B));
INV_X1 FE_OFC83_g2176B (.ZN(FE_OFN83_g2176B),.A(FE_OFN81_g2176B));
INV_X1 FE_OFC82_g2176B (.ZN(FE_OFN82_g2176B),.A(FE_OFN81_g2176B));
INV_X1 FE_OFC81_g2176B (.ZN(FE_OFN81_g2176B),.A(g2176B));
BUF_X3 FE_OFC80_g2175B (.Z(FE_OFN80_g2175B),.A(g2175B));
INV_X1 FE_OFC79_g8700B (.ZN(FE_OFN79_g8700B),.A(g9097B));
BUF_X3 FE_OFC76_g8700B (.Z(FE_OFN76_g8700B),.A(g8700B));
BUF_X3 FE_OFC73_g8858B (.Z(FE_OFN73_g8858B),.A(g8858B));
BUF_X3 FE_OFC72_g9292B (.Z(FE_OFN72_g9292B),.A(FE_OFN71_g9292B));
BUF_X3 FE_OFC71_g9292B (.Z(FE_OFN71_g9292B),.A(g9292B));
BUF_X3 FE_OFC70_g9490B (.Z(FE_OFN70_g9490B),.A(g9490B));
BUF_X3 FE_OFC69_g9392B (.Z(FE_OFN69_g9392B),.A(FE_OFN68_g9392B));
BUF_X3 FE_OFC68_g9392B (.Z(FE_OFN68_g9392B),.A(g9392B));
BUF_X3 FE_OFC67_g9367B (.Z(FE_OFN67_g9367B),.A(g9367B));
BUF_X3 FE_OFC64_g9536B (.Z(FE_OFN64_g9536B),.A(g9536B));
BUF_X3 FE_OFC63_g9474B (.Z(FE_OFN63_g9474B),.A(g9474B));
BUF_X3 FE_OFC62_g9274B (.Z(FE_OFN62_g9274B),.A(g9274B));
BUF_X3 FE_OFC61_g9624B (.Z(FE_OFN61_g9624B),.A(FE_OFN60_g9624B));
BUF_X3 FE_OFC60_g9624B (.Z(FE_OFN60_g9624B),.A(g9624B));
INV_X1 FE_OFC59_g9432B (.ZN(FE_OFN59_g9432B),.A(FE_OFN57_g9432B));
INV_X1 FE_OFC57_g9432B (.ZN(FE_OFN57_g9432B),.A(g9432B));
BUF_X3 FE_OFC56_g9052B (.Z(FE_OFN56_g9052B),.A(FE_OFN54_g9052B));
BUF_X3 FE_OFC54_g9052B (.Z(FE_OFN54_g9052B),.A(g9052B));
BUF_X3 FE_OFC53_g9173B (.Z(FE_OFN53_g9173B),.A(FE_OFN52_g9173B));
BUF_X3 FE_OFC52_g9173B (.Z(FE_OFN52_g9173B),.A(g9173B));
BUF_X3 FE_OFC51_g9111B (.Z(FE_OFN51_g9111B),.A(g9111B));
BUF_X3 FE_OFC50_g9030B (.Z(FE_OFN50_g9030B),.A(FE_OFN49_g9030B));
BUF_X3 FE_OFC49_g9030B (.Z(FE_OFN49_g9030B),.A(g9030B));
BUF_X3 FE_OFC48_g9151B (.Z(FE_OFN48_g9151B),.A(FE_OFN47_g9151B));
BUF_X3 FE_OFC47_g9151B (.Z(FE_OFN47_g9151B),.A(g9151B));
BUF_X3 FE_OFC46_g9125B (.Z(FE_OFN46_g9125B),.A(FE_OFN45_g9125B));
BUF_X3 FE_OFC45_g9125B (.Z(FE_OFN45_g9125B),.A(FE_OFN44_g9125B));
BUF_X3 FE_OFC44_g9125B (.Z(FE_OFN44_g9125B),.A(g9125B));
BUF_X3 FE_OFC42_g9205B (.Z(FE_OFN42_g9205B),.A(g9205B));
BUF_X3 FE_OFC40_g9240B (.Z(FE_OFN40_g9240B),.A(g9240B));
BUF_X3 FE_OFC39_g9223B (.Z(FE_OFN39_g9223B),.A(g9223B));
BUF_X3 FE_OFC35_g9785B (.Z(FE_OFN35_g9785B),.A(FE_OFN34_g9785B));
BUF_X3 FE_OFC34_g9785B (.Z(FE_OFN34_g9785B),.A(g9785B));
BUF_X3 FE_OFC33_g9454B (.Z(FE_OFN33_g9454B),.A(FE_OFN32_g9454B));
BUF_X3 FE_OFC32_g9454B (.Z(FE_OFN32_g9454B),.A(g9454B));
BUF_X3 FE_OFC27_g11519B (.Z(FE_OFN27_g11519B),.A(g11519B));
BUF_X3 FE_OFC21_g10702B (.Z(FE_OFN21_g10702B),.A(FE_OFN20_g10702B));
BUF_X3 FE_OFC20_g10702B (.Z(FE_OFN20_g10702B),.A(FE_OFN18_g10702B));
BUF_X3 FE_OFC18_g10702B (.Z(FE_OFN18_g10702B),.A(FE_OFN13_g10702B));
INV_X1 FE_OFC17_g10702B (.ZN(FE_OFN17_g10702B),.A(FE_OFN15_g10702B));
INV_X1 FE_OFC15_g10702B (.ZN(FE_OFN15_g10702B),.A(FE_OFN14_g10702B));
BUF_X3 FE_OFC14_g10702B (.Z(FE_OFN14_g10702B),.A(FE_OFN9_g10702B));
INV_X1 FE_OFC13_g10702B (.ZN(FE_OFN13_g10702B),.A(FE_OFN10_g10702B));
INV_X1 FE_OFC10_g10702B (.ZN(FE_OFN10_g10702B),.A(FE_OFN9_g10702B));
BUF_X3 FE_OFC9_g10702B (.Z(FE_OFN9_g10702B),.A(FE_OFN8_g10702B));
BUF_X3 FE_OFC8_g10702B (.Z(FE_OFN8_g10702B),.A(FE_OFN7_g10702B));
BUF_X3 FE_OFC7_g10702B (.Z(FE_OFN7_g10702B),.A(g10702B));
BUF_X3 FE_OFC4_g10950B (.Z(FE_OFN4_g10950B),.A(FE_OFN3_g10950B));
INV_X1 FE_OFC3_g10950B (.ZN(FE_OFN3_g10950B),.A(FE_OFN0_g10950B));
INV_X1 FE_OFC0_g10950B (.ZN(FE_OFN0_g10950B),.A(g10950B));
INV_X1 U_g2299B (.ZN(g2299B),.A(g1707B));
INV_X1 U_g9291B (.ZN(g9291B),.A(FE_OFN79_g8700B));
INV_X4 U_I7048B (.ZN(I7048B),.A(g2807B));
INV_X1 U_g1981B (.ZN(g1981B),.A(g650B));
INV_X1 U_g3982B (.ZN(g3982B),.A(g2118B));
INV_X1 U_g3629B (.ZN(g3629B),.A(FE_OFN266_g18B));
INV_X1 U_g6842B (.ZN(g6842B),.A(I9769B));
INV_X1 U_g8617B (.ZN(g8617B),.A(g8465B));
INV_X1 U_g2078B (.ZN(g2078B),.A(g135B));
INV_X1 U_g2340B (.ZN(g2340B),.A(g1918B));
INV_X1 U_g7684B (.ZN(g7684B),.A(FE_OFN83_g2176B));
INV_X1 U_g3800B (.ZN(g3800B),.A(FE_OFN250_g471B));
INV_X1 U_g6941B (.ZN(g6941B),.A(FE_OFN88_g2178B));
INV_X1 U_g2435B (.ZN(g2435B),.A(g201B));
INV_X4 U_g4010B (.ZN(g4010B),.A(g3744B));
INV_X1 U_g2082B (.ZN(g2082B),.A(g1371B));
INV_X1 U_g5519B (.ZN(g5519B),.A(g4811B));
INV_X1 U_g10668B (.ZN(g10668B),.A(g10563B));
INV_X1 U_g4172B (.ZN(g4172B),.A(g2057B));
INV_X1 U_g8709B (.ZN(g8709B),.A(g8451B));
INV_X1 U_g2214B (.ZN(g2214B),.A(g115B));
INV_X1 U_I7847B (.ZN(I7847B),.A(g3435B));
INV_X1 U_g8340B (.ZN(g8340B),.A(I13400B));
INV_X1 U_g4566B (.ZN(g4566B),.A(g3753B));
INV_X1 U_g3348B (.ZN(g3348B),.A(FE_OFN267_g109B));
INV_X1 U_I15968B (.ZN(I15968B),.A(g10408B));
INV_X1 U_g11060B (.ZN(g11060B),.A(g10937B));
INV_X1 U_I15855B (.ZN(I15855B),.A(g10336B));
INV_X1 U_g6270B (.ZN(g6270B),.A(I9383B));
INV_X1 U_g10679B (.ZN(g10679B),.A(g10584B));
INV_X1 U_g1968B (.ZN(g1968B),.A(g369B));
INV_X1 U_g5659B (.ZN(g5659B),.A(I7771B));
INV_X1 U_I15503B (.ZN(I15503B),.A(g9995B));
INV_X1 U_g8110B (.ZN(g8110B),.A(g7996B));
INV_X1 U_g2556B (.ZN(g2556B),.A(g186B));
INV_X1 U_I7817B (.ZN(I7817B),.A(g3399B));
INV_X1 U_g2222B (.ZN(g2222B),.A(g158B));
INV_X1 U_I13373B (.ZN(I13373B),.A(g8226B));
INV_X1 U_g4202B (.ZN(g4202B),.A(I5430B));
INV_X1 U_I9880B (.ZN(I9880B),.A(g5405B));
INV_X1 U_g4094B (.ZN(g4094B),.A(g2744B));
INV_X1 U_g4567B (.ZN(g4567B),.A(g3374B));
INV_X1 U_I14312B (.ZN(I14312B),.A(g8814B));
INV_X1 U_g11111B (.ZN(g11111B),.A(g10702B));
INV_X1 U_g4776B (.ZN(g4776B),.A(FE_OFN344_g3586B));
INV_X1 U_I15986B (.ZN(I15986B),.A(g10417B));
INV_X1 U_g2237B (.ZN(g2237B),.A(g713B));
INV_X1 U_g7897B (.ZN(g7897B),.A(g7712B));
INV_X1 U_g3121B (.ZN(g3121B),.A(FE_OFN352_g109B));
INV_X1 U_g5420B (.ZN(g5420B),.A(g4300B));
INV_X1 U_g10455B (.ZN(g10455B),.A(I15956B));
INV_X1 U_g2557B (.ZN(g2557B),.A(g1840B));
INV_X1 U_g9097B (.ZN(g9097B),.A(g8700B));
INV_X1 U_g3938B (.ZN(g3938B),.A(g2299B));
INV_X1 U_g8563B (.ZN(g8563B),.A(I7829B));
INV_X1 U_g6259B (.ZN(g6259B),.A(g2175B));
INV_X1 U_g4179B (.ZN(g4179B),.A(g1992B));
INV_X1 U_g7682B (.ZN(g7682B),.A(FE_OFN83_g2176B));
INV_X1 U_g4379B (.ZN(g4379B),.A(g3698B));
INV_X1 U_I4917B (.ZN(I4917B),.A(g584B));
INV_X1 U_g2254B (.ZN(g2254B),.A(g131B));
INV_X1 U_g4289B (.ZN(g4289B),.A(FE_OFN298_g3015B));
INV_X1 U_g4777B (.ZN(g4777B),.A(g3992B));
INV_X1 U_g8089B (.ZN(g8089B),.A(g7934B));
INV_X1 U_g2438B (.ZN(g2438B),.A(g243B));
INV_X1 U_g4271B (.ZN(g4271B),.A(g2024B));
INV_X1 U_g7045B (.ZN(g7045B),.A(g6003B));
INV_X1 U_I5424B (.ZN(I5424B),.A(g910B));
INV_X1 U_g2212B (.ZN(g2212B),.A(g686B));
INV_X1 U_g3141B (.ZN(g3141B),.A(g2563B));
INV_X1 U_g3710B (.ZN(g3710B),.A(g3215B));
INV_X1 U_g7920B (.ZN(g7920B),.A(g7516B));
INV_X1 U_g2229B (.ZN(g2229B),.A(g162B));
INV_X1 U_I15157B (.ZN(I15157B),.A(g9931B));
INV_X1 U_g11157B (.ZN(g11157B),.A(FE_OFN3_g10950B));
INV_X1 U_g4209B (.ZN(g4209B),.A(I5002B));
INV_X1 U_I9279B (.ZN(I9279B),.A(g91B));
INV_X1 U_I5044B (.ZN(I5044B),.A(g1182B));
INV_X1 U_I15287B (.ZN(I15287B),.A(g9968B));
INV_X1 U_g2249B (.ZN(g2249B),.A(g127B));
INV_X1 U_g11596B (.ZN(g11596B),.A(g11580B));
INV_X1 U_g11243B (.ZN(g11243B),.A(FE_OFN8_g10702B));
INV_X1 U_g6266B (.ZN(g6266B),.A(g2208B));
INV_X1 U_g8062B (.ZN(g8062B),.A(I4783B));
INV_X1 U_I5414B (.ZN(I5414B),.A(g904B));
INV_X1 U_g3628B (.ZN(g3628B),.A(g3111B));
INV_X1 U_g6255B (.ZN(g6255B),.A(I9237B));
INV_X1 U_g4175B (.ZN(g4175B),.A(g1988B));
INV_X1 U_g6081B (.ZN(g6081B),.A(g4977B));
INV_X1 U_g7910B (.ZN(g7910B),.A(g7460B));
INV_X1 U_g4285B (.ZN(g4285B),.A(g3688B));
INV_X1 U_g6354B (.ZN(g6354B),.A(g5867B));
INV_X1 U_g2031B (.ZN(g2031B),.A(g1690B));
INV_X1 U_g8085B (.ZN(g8085B),.A(g7932B));
INV_X1 U_g2176B (.ZN(g2176B),.A(g82B));
INV_X1 U_g7883B (.ZN(g7883B),.A(g7246B));
INV_X1 U_g4737B (.ZN(g4737B),.A(g3440B));
INV_X1 U_I13351B (.ZN(I13351B),.A(g8214B));
INV_X1 U_g6267B (.ZN(g6267B),.A(I9326B));
INV_X1 U_g3440B (.ZN(g3440B),.A(g3041B));
INV_X1 U_g2610B (.ZN(g2610B),.A(I4917B));
INV_X1 U_g4205B (.ZN(g4205B),.A(I4992B));
INV_X1 U_g10883B (.ZN(g10883B),.A(g10809B));
INV_X1 U_g5521B (.ZN(g5521B),.A(FE_OFN221_g3440B));
INV_X1 U_I6260B (.ZN(I6260B),.A(g1696B));
INV_X1 U_I9311B (.ZN(I9311B),.A(g103B));
INV_X1 U_I5579B (.ZN(I5579B),.A(g1197B));
INV_X1 U_g10439B (.ZN(g10439B),.A(g10334B));
INV_X1 U_g5878B (.ZN(g5878B),.A(g5309B));
INV_X1 U_g6932B (.ZN(g6932B),.A(I7829B));
INV_X1 U_g4273B (.ZN(g4273B),.A(FE_OFN133_g3015B));
INV_X1 U_g5658B (.ZN(g5658B),.A(I7752B));
INV_X1 U_g7467B (.ZN(g7467B),.A(FE_OFN84_g2176B));
INV_X1 U_g1990B (.ZN(g1990B),.A(g774B));
INV_X1 U_I13436B (.ZN(I13436B),.A(g8187B));
INV_X1 U_g2399B (.ZN(g2399B),.A(g605B));
INV_X1 U_g8980B (.ZN(g8980B),.A(I14306B));
INV_X1 U_g6716B (.ZN(g6716B),.A(FE_OFN115_g4807B));
INV_X1 U_g7685B (.ZN(g7685B),.A(FE_OFN87_g2176B));
INV_X1 U_g8849B (.ZN(g8849B),.A(g8745B));
INV_X1 U_I7840B (.ZN(I7840B),.A(g3431B));
INV_X1 U_g10852B (.ZN(g10852B),.A(g10739B));
INV_X1 U_g7562B (.ZN(g7562B),.A(FE_OFN91_g2172B));
INV_X1 U_g6258B (.ZN(g6258B),.A(g2172B));
INV_X1 U_g4178B (.ZN(g4178B),.A(g1991B));
INV_X4 U_g4679B (.ZN(g4679B),.A(FE_OFN293_g3015B));
INV_X1 U_g3776B (.ZN(g3776B),.A(g2579B));
INV_X1 U_g2008B (.ZN(g2008B),.A(g971B));
INV_X1 U_g6274B (.ZN(g6274B),.A(I9293B));
INV_X1 U_g2336B (.ZN(g2336B),.A(g1900B));
INV_X1 U_g3521B (.ZN(g3521B),.A(FE_OFN359_g18B));
INV_X1 U_g6280B (.ZN(g6280B),.A(g2253B));
INV_X1 U_I6962B (.ZN(I6962B),.A(g2791B));
INV_X1 U_g2230B (.ZN(g2230B),.A(g704B));
INV_X1 U_g4437B (.ZN(g4437B),.A(FE_OFN235_g2024B));
INV_X1 U_g4208B (.ZN(g4208B),.A(I5588B));
INV_X1 U_g7505B (.ZN(g7505B),.A(FE_OFN87_g2176B));
INV_X1 U_I15974B (.ZN(I15974B),.A(g10411B));
INV_X1 U_g2550B (.ZN(g2550B),.A(g1834B));
INV_X1 U_g10400B (.ZN(g10400B),.A(g10348B));
INV_X1 U_I9282B (.ZN(I9282B),.A(g101B));
INV_X1 U_I5584B (.ZN(I5584B),.A(g1200B));
INV_X4 U_g9490B (.ZN(g9490B),.A(g9324B));
INV_X1 U_g2395B (.ZN(g2395B),.A(g231B));
INV_X1 U_g8465B (.ZN(g8465B),.A(g8289B));
INV_X1 U_g6403B (.ZN(g6403B),.A(g5013B));
INV_X1 U_I15510B (.ZN(I15510B),.A(g10013B));
INV_X1 U_g2248B (.ZN(g2248B),.A(g99B));
INV_X1 U_g3744B (.ZN(g3744B),.A(FE_OFN269_g109B));
INV_X1 U_I4883B (.ZN(I4883B),.A(g581B));
INV_X1 U_g7688B (.ZN(g7688B),.A(FE_OFN83_g2176B));
INV_X1 U_g2481B (.ZN(g2481B),.A(g882B));
INV_X1 U_g10683B (.ZN(g10683B),.A(g10385B));
INV_X1 U_I5070B (.ZN(I5070B),.A(g1194B));
INV_X1 U_g4888B (.ZN(g4888B),.A(I5101B));
INV_X1 U_g4171B (.ZN(g4171B),.A(I6962B));
INV_X1 U_g4787B (.ZN(g4787B),.A(g3423B));
INV_X1 U_g6447B (.ZN(g6447B),.A(FE_OFN218_g5557B));
INV_X1 U_g3092B (.ZN(g3092B),.A(g639B));
INV_X1 U_g4281B (.ZN(g4281B),.A(g3586B));
INV_X1 U_g5613B (.ZN(g5613B),.A(FE_OFN131_g3015B));
INV_X1 U_g8255B (.ZN(g8255B),.A(g7986B));
INV_X1 U_g8081B (.ZN(g8081B),.A(g8000B));
INV_X1 U_I5406B (.ZN(I5406B),.A(g898B));
INV_X1 U_I4780B (.ZN(I4780B),.A(g872B));
INV_X1 U_g10584B (.ZN(g10584B),.A(g10522B));
INV_X1 U_g6272B (.ZN(g6272B),.A(I9268B));
INV_X1 U_g8783B (.ZN(g8783B),.A(g8746B));
INV_X1 U_g8979B (.ZN(g8979B),.A(I14303B));
INV_X1 U_g4201B (.ZN(g4201B),.A(I5427B));
INV_X1 U_I5445B (.ZN(I5445B),.A(g922B));
INV_X1 U_g4449B (.ZN(g4449B),.A(g4144B));
INV_X1 U_g7696B (.ZN(g7696B),.A(FE_OFN86_g2176B));
INV_X1 U_g8828B (.ZN(g8828B),.A(g8744B));
INV_X1 U_g2677B (.ZN(g2677B),.A(g2034B));
INV_X1 U_g10361B (.ZN(g10361B),.A(g10268B));
INV_X1 U_g3737B (.ZN(g3737B),.A(g2506B));
INV_X1 U_I9332B (.ZN(I9332B),.A(g104B));
INV_X1 U_g9525B (.ZN(g9525B),.A(g9257B));
INV_X1 U_g2198B (.ZN(g2198B),.A(g668B));
INV_X1 U_I7771B (.ZN(I7771B),.A(g3418B));
INV_X1 U_g3523B (.ZN(g3523B),.A(g1845B));
INV_X1 U_g2241B (.ZN(g2241B),.A(g722B));
INV_X1 U_g7681B (.ZN(g7681B),.A(FE_OFN87_g2176B));
INV_X1 U_g7697B (.ZN(g7697B),.A(g7101B));
INV_X1 U_g7914B (.ZN(g7914B),.A(g7651B));
INV_X1 U_g8349B (.ZN(g8349B),.A(I13427B));
INV_X1 U_g6260B (.ZN(g6260B),.A(g2178B));
INV_X1 U_I14319B (.ZN(I14319B),.A(g8816B));
INV_X1 U_g10463B (.ZN(g10463B),.A(I15980B));
INV_X1 U_I5388B (.ZN(I5388B),.A(g889B));
INV_X1 U_g2211B (.ZN(g2211B),.A(g153B));
INV_X1 U_g6279B (.ZN(g6279B),.A(g2248B));
INV_X1 U_g3983B (.ZN(g3983B),.A(g3222B));
INV_X1 U_I5430B (.ZN(I5430B),.A(g916B));
INV_X4 U_g4678B (.ZN(g4678B),.A(g3546B));
INV_X1 U_g3543B (.ZN(g3543B),.A(g3101B));
INV_X1 U_g9507B (.ZN(g9507B),.A(g9268B));
INV_X1 U_g10421B (.ZN(g10421B),.A(g10331B));
INV_X1 U_g8352B (.ZN(g8352B),.A(I13436B));
INV_X1 U_g7460B (.ZN(g7460B),.A(FE_OFN85_g2176B));
INV_X1 U_g2083B (.ZN(g2083B),.A(g139B));
INV_X1 U_I6360B (.ZN(I6360B),.A(g1713B));
INV_X1 U_I4992B (.ZN(I4992B),.A(g1170B));
INV_X1 U_I16982B (.ZN(I16982B),.A(g10629B));
INV_X1 U_g8599B (.ZN(g8599B),.A(g8546B));
INV_X1 U_g6253B (.ZN(g6253B),.A(I9479B));
INV_X1 U_g2061B (.ZN(g2061B),.A(g1828B));
INV_X1 U_g2187B (.ZN(g2187B),.A(g746B));
INV_X1 U_g4173B (.ZN(g4173B),.A(g1984B));
INV_X1 U_g8984B (.ZN(g8984B),.A(I14319B));
INV_X1 U_g2446B (.ZN(g2446B),.A(g1400B));
INV_X1 U_g11575B (.ZN(g11575B),.A(g11561B));
INV_X1 U_g2345B (.ZN(g2345B),.A(g1936B));
INV_X1 U_g8106B (.ZN(g8106B),.A(g7950B));
INV_X1 U_g6586B (.ZN(g6586B),.A(FE_OFN118_g4807B));
INV_X1 U_g8061B (.ZN(g8061B),.A(I4780B));
INV_X1 U_g5808B (.ZN(g5808B),.A(g85B));
INV_X1 U_I5418B (.ZN(I5418B),.A(g907B));
INV_X1 U_g4203B (.ZN(g4203B),.A(I5441B));
INV_X1 U_g2016B (.ZN(g2016B),.A(g1361B));
INV_X1 U_I16252B (.ZN(I16252B),.A(g10515B));
INV_X1 U_I9273B (.ZN(I9273B),.A(g47B));
INV_X1 U_g2251B (.ZN(g2251B),.A(g731B));
INV_X1 U_g2047B (.ZN(g2047B),.A(g1857B));
INV_X1 U_g10927B (.ZN(g10927B),.A(FE_OFN17_g10702B));
INV_X1 U_g6275B (.ZN(g6275B),.A(I9308B));
INV_X1 U_g4216B (.ZN(g4216B),.A(I5070B));
INV_X1 U_g8858B (.ZN(g8858B),.A(g8743B));
INV_X1 U_g4671B (.ZN(g4671B),.A(g3354B));
INV_X1 U_g8115B (.ZN(g8115B),.A(g7953B));
INV_X1 U_g2612B (.ZN(g2612B),.A(I4948B));
INV_X1 U_g2017B (.ZN(g2017B),.A(g1218B));
INV_X1 U_g6284B (.ZN(g6284B),.A(I9332B));
INV_X1 U_g7683B (.ZN(g7683B),.A(FE_OFN87_g2176B));
INV_X1 U_I5101B (.ZN(I5101B),.A(g1960B));
INV_X1 U_g2328B (.ZN(g2328B),.A(g1882B));
INV_X1 U_g2542B (.ZN(g2542B),.A(g1868B));
INV_X1 U_g2330B (.ZN(g2330B),.A(g1891B));
INV_X1 U_g7949B (.ZN(g7949B),.A(FE_OFN211_g7246B));
INV_X1 U_I5041B (.ZN(I5041B),.A(g1179B));
INV_X1 U_g1992B (.ZN(g1992B),.A(g782B));
INV_X1 U_g8978B (.ZN(g8978B),.A(I14299B));
INV_X1 U_I5441B (.ZN(I5441B),.A(g919B));
INV_X1 U_g4365B (.ZN(g4365B),.A(g3880B));
INV_X1 U_g8982B (.ZN(g8982B),.A(I14312B));
INV_X1 U_g8234B (.ZN(g8234B),.A(FE_OFN198_g7697B));
INV_X1 U_g8328B (.ZN(g8328B),.A(I13364B));
INV_X1 U_g4196B (.ZN(g4196B),.A(I5245B));
INV_X1 U_g2456B (.ZN(g2456B),.A(g1397B));
INV_X1 U_g7919B (.ZN(g7919B),.A(g7512B));
INV_X1 U_g5105B (.ZN(g5105B),.A(I4783B));
INV_X1 U_g1976B (.ZN(g1976B),.A(g643B));
INV_X1 U_g7952B (.ZN(g7952B),.A(FE_OFN210_g7246B));
INV_X1 U_I4820B (.ZN(I4820B),.A(g865B));
INV_X1 U_g2355B (.ZN(g2355B),.A(I5435B));
INV_X1 U_I14315B (.ZN(I14315B),.A(g8815B));
INV_X1 U_g4467B (.ZN(g4467B),.A(g3829B));
INV_X1 U_g4290B (.ZN(g4290B),.A(FE_OFN102_g3586B));
INV_X1 U_g7527B (.ZN(g7527B),.A(FE_OFN85_g2176B));
INV_X1 U_I9265B (.ZN(I9265B),.A(g46B));
INV_X1 U_g8056B (.ZN(g8056B),.A(g7671B));
INV_X1 U_g4181B (.ZN(g4181B),.A(g2449B));
INV_X1 U_g4381B (.ZN(g4381B),.A(FE_OFN296_g3914B));
INV_X1 U_g2118B (.ZN(g2118B),.A(g1854B));
INV_X1 U_I6273B (.ZN(I6273B),.A(FE_OFN363_I5565B));
INV_X1 U_g10629B (.ZN(g10629B),.A(g10583B));
INV_X1 U_g4197B (.ZN(g4197B),.A(I5410B));
INV_X1 U_g2652B (.ZN(g2652B),.A(g2008B));
INV_X1 U_g2057B (.ZN(g2057B),.A(g754B));
INV_X1 U_g10628B (.ZN(g10628B),.A(I16252B));
INV_X1 U_g3539B (.ZN(g3539B),.A(g3015B));
INV_X1 U_g4263B (.ZN(g4263B),.A(FE_OFN103_g3586B));
INV_X1 U_I9296B (.ZN(I9296B),.A(g102B));
INV_X1 U_I13323B (.ZN(I13323B),.A(g8203B));
INV_X1 U_g2549B (.ZN(g2549B),.A(g1386B));
INV_X1 U_g6278B (.ZN(g6278B),.A(I9371B));
INV_X1 U_g5261B (.ZN(g5261B),.A(g4640B));
INV_X1 U_g3419B (.ZN(g3419B),.A(g3104B));
INV_X1 U_I7829B (.ZN(I7829B),.A(g3425B));
INV_X1 U_g7516B (.ZN(g7516B),.A(FE_OFN82_g2176B));
INV_X1 U_g6282B (.ZN(g6282B),.A(I9296B));
INV_X1 U_g9802B (.ZN(g9802B),.A(g9490B));
INV_X1 U_g8318B (.ZN(g8318B),.A(I13338B));
INV_X1 U_g3086B (.ZN(g3086B),.A(g2276B));
INV_X1 U_g2253B (.ZN(g2253B),.A(g100B));
INV_X1 U_I9371B (.ZN(I9371B),.A(g96B));
INV_X1 U_I5383B (.ZN(I5383B),.A(g886B));
INV_X1 U_g2606B (.ZN(g2606B),.A(I4876B));
INV_X1 U_I5588B (.ZN(I5588B),.A(g1203B));
INV_X1 U_g7907B (.ZN(g7907B),.A(g7664B));
INV_X1 U_g4673B (.ZN(g4673B),.A(FE_OFN348_g3015B));
INV_X1 U_g2570B (.ZN(g2570B),.A(g207B));
INV_X1 U_g7915B (.ZN(g7915B),.A(g7473B));
INV_X1 U_g10377B (.ZN(g10377B),.A(I15855B));
INV_X1 U_g6264B (.ZN(g6264B),.A(g2176B));
INV_X1 U_g2607B (.ZN(g2607B),.A(I4883B));
INV_X1 U_g2506B (.ZN(g2506B),.A(g636B));
INV_X1 U_I16717B (.ZN(I16717B),.A(g10779B));
INV_X1 U_g3491B (.ZN(g3491B),.A(g1107B));
INV_X1 U_I7852B (.ZN(I7852B),.A(g3438B));
INV_X1 U_g2275B (.ZN(g2275B),.A(g757B));
INV_X1 U_g3007B (.ZN(g3007B),.A(I6240B));
INV_X1 U_g2374B (.ZN(g2374B),.A(g591B));
INV_X1 U_I9268B (.ZN(I9268B),.A(g90B));
INV_X1 U_g9424B (.ZN(g9424B),.A(g9291B));
INV_X1 U_g6271B (.ZN(g6271B),.A(I9259B));
INV_X1 U_g3793B (.ZN(g3793B),.A(FE_OFN248_g466B));
INV_X1 U_I7825B (.ZN(I7825B),.A(g3414B));
INV_X1 U_g2420B (.ZN(g2420B),.A(g237B));
INV_X1 U_g3664B (.ZN(g3664B),.A(g3209B));
INV_X1 U_g5509B (.ZN(g5509B),.A(g4739B));
INV_X1 U_g8985B (.ZN(g8985B),.A(I14326B));
INV_X1 U_g4608B (.ZN(g4608B),.A(FE_OFN141_g3829B));
INV_X1 U_g5816B (.ZN(g5816B),.A(g1810B));
INV_X1 U_I5060B (.ZN(I5060B),.A(g1191B));
INV_X1 U_I14306B (.ZN(I14306B),.A(g8812B));
INV_X1 U_g9961B (.ZN(g9961B),.A(I15157B));
INV_X1 U_g7438B (.ZN(g7438B),.A(FE_OFN195_g6488B));
INV_X1 U_g8100B (.ZN(g8100B),.A(g7947B));
INV_X1 U_g5101B (.ZN(g5101B),.A(I4780B));
INV_X1 U_g7918B (.ZN(g7918B),.A(g7505B));
INV_X1 U_g6262B (.ZN(g6262B),.A(I9273B));
INV_X1 U_g2648B (.ZN(g2648B),.A(I4820B));
INV_X1 U_g2410B (.ZN(g2410B),.A(g1453B));
INV_X1 U_g8323B (.ZN(g8323B),.A(I13351B));
INV_X1 U_I5053B (.ZN(I5053B),.A(g1188B));
INV_X1 U_g6285B (.ZN(g6285B),.A(I9352B));
INV_X1 U_g2172B (.ZN(g2172B),.A(g43B));
INV_X1 U_I13364B (.ZN(I13364B),.A(g8221B));
INV_X1 U_g2343B (.ZN(g2343B),.A(g1927B));
INV_X1 U_g4210B (.ZN(g4210B),.A(I5020B));
INV_X1 U_I4876B (.ZN(I4876B),.A(g580B));
INV_X1 U_g8566B (.ZN(g8566B),.A(I7852B));
INV_X1 U_g2202B (.ZN(g2202B),.A(g148B));
INV_X1 U_g6926B (.ZN(g6926B),.A(I7825B));
INV_X1 U_g8548B (.ZN(g8548B),.A(g8390B));
INV_X1 U_g2518B (.ZN(g2518B),.A(g590B));
INV_X1 U_g6273B (.ZN(g6273B),.A(I9279B));
INV_X1 U_g10801B (.ZN(g10801B),.A(I16507B));
INV_X1 U_g4739B (.ZN(g4739B),.A(g4117B));
INV_X1 U_g6269B (.ZN(g6269B),.A(I9368B));
INV_X1 U_g8313B (.ZN(g8313B),.A(I13323B));
INV_X1 U_I9308B (.ZN(I9308B),.A(g93B));
INV_X1 U_g4294B (.ZN(g4294B),.A(g3664B));
INV_X1 U_g3723B (.ZN(g3723B),.A(g3071B));
INV_X1 U_g10457B (.ZN(g10457B),.A(I15962B));
INV_X1 U_g8094B (.ZN(g8094B),.A(g7987B));
INV_X1 U_g2050B (.ZN(g2050B),.A(g1861B));
INV_X1 U_g7473B (.ZN(g7473B),.A(FE_OFN87_g2176B));
INV_X1 U_g2777B (.ZN(g2777B),.A(FE_OFN224_g2276B));
INV_X1 U_g2271B (.ZN(g2271B),.A(g877B));
INV_X1 U_g2611B (.ZN(g2611B),.A(I4935B));
INV_X1 U_g3368B (.ZN(g3368B),.A(g2459B));
INV_X1 U_g1987B (.ZN(g1987B),.A(g762B));
INV_X4 U_I8869B (.ZN(I8869B),.A(g4421B));
INV_X1 U_I9290B (.ZN(I9290B),.A(FE_OFN277_g48B));
INV_X1 U_I4948B (.ZN(I4948B),.A(g586B));
INV_X1 U_g8271B (.ZN(g8271B),.A(g1810B));
INV_X1 U_g1991B (.ZN(g1991B),.A(g778B));
INV_X1 U_g11199B (.ZN(g11199B),.A(FE_OFN21_g10702B));
INV_X1 U_g8981B (.ZN(g8981B),.A(I14309B));
INV_X1 U_I15365B (.ZN(I15365B),.A(g10025B));
INV_X1 U_g7852B (.ZN(g7852B),.A(FE_OFN209_g6863B));
INV_X1 U_g7923B (.ZN(g7923B),.A(g7527B));
INV_X1 U_g10431B (.ZN(g10431B),.A(g10328B));
INV_X1 U_g6265B (.ZN(g6265B),.A(I9276B));
INV_X1 U_g4782B (.ZN(g4782B),.A(g4089B));
INV_X1 U_g4292B (.ZN(g4292B),.A(FE_OFN136_g3863B));
INV_X1 U_g3760B (.ZN(g3760B),.A(g3003B));
INV_X1 U_I5435B (.ZN(I5435B),.A(g18B));
INV_X1 U_g5117B (.ZN(g5117B),.A(FE_OFN144_g4682B));
INV_X4 U_g2175B (.ZN(g2175B),.A(g44B));
INV_X1 U_I9368B (.ZN(I9368B),.A(g87B));
INV_X4 U_g2024B (.ZN(g2024B),.A(g1718B));
INV_X1 U_g6281B (.ZN(g6281B),.A(I9282B));
INV_X1 U_g3327B (.ZN(g3327B),.A(g23B));
INV_X4 U_g2424B (.ZN(g2424B),.A(FE_OFN241_g1690B));
INV_X1 U_I5002B (.ZN(I5002B),.A(g1173B));
INV_X1 U_g7550B (.ZN(g7550B),.A(FE_OFN96_g2169B));
INV_X1 U_g2077B (.ZN(g2077B),.A(g219B));
INV_X1 U_g3103B (.ZN(g3103B),.A(g1212B));
INV_X1 U_g7913B (.ZN(g7913B),.A(g7467B));
INV_X1 U_g6109B (.ZN(g6109B),.A(g48B));
INV_X1 U_g6449B (.ZN(g6449B),.A(g5557B));
INV_X1 U_g2273B (.ZN(g2273B),.A(g881B));
INV_X1 U_g7692B (.ZN(g7692B),.A(g2176B));
INV_X1 U_g7497B (.ZN(g7497B),.A(FE_OFN85_g2176B));
INV_X1 U_g2444B (.ZN(g2444B),.A(g876B));
INV_X1 U_g8099B (.ZN(g8099B),.A(g7990B));
INV_X1 U_I9326B (.ZN(I9326B),.A(FE_OFN271_g85B));
INV_X1 U_g6268B (.ZN(g6268B),.A(I9346B));
INV_X1 U_g10676B (.ZN(g10676B),.A(g10570B));
INV_X1 U_g1993B (.ZN(g1993B),.A(g786B));
INV_X1 U_I9383B (.ZN(I9383B),.A(g88B));
INV_X1 U_g8983B (.ZN(g8983B),.A(I14315B));
INV_X1 U_I5254B (.ZN(I5254B),.A(g1700B));
INV_X1 U_I14303B (.ZN(I14303B),.A(g8811B));
INV_X1 U_g2178B (.ZN(g2178B),.A(g45B));
INV_X1 U_I4900B (.ZN(I4900B),.A(g583B));
INV_X1 U_g3060B (.ZN(g3060B),.A(FE_OFN245_g1690B));
INV_X1 U_g4214B (.ZN(g4214B),.A(I5053B));
INV_X1 U_I9346B (.ZN(I9346B),.A(g86B));
INV_X1 U_g2382B (.ZN(g2382B),.A(g599B));
INV_X1 U_g3784B (.ZN(g3784B),.A(FE_OFN254_g461B));
INV_X1 U_I17413B (.ZN(I17413B),.A(g11425B));
INV_X1 U_g7677B (.ZN(g7677B),.A(FE_OFN85_g2176B));
INV_X4 U_g4002B (.ZN(g4002B),.A(FE_OFN155_g3121B));
INV_X1 U_g3479B (.ZN(g3479B),.A(g1101B));
INV_X1 U_g11489B (.ZN(g11489B),.A(I17413B));
INV_X1 U_g6131B (.ZN(g6131B),.A(g5548B));
INV_X1 U_g3390B (.ZN(g3390B),.A(g2045B));
INV_X1 U_g5627B (.ZN(g5627B),.A(FE_OFN132_g3015B));
INV_X1 U_g3501B (.ZN(g3501B),.A(FE_OFN240_g1110B));
INV_X1 U_g8335B (.ZN(g8335B),.A(I13385B));
INV_X1 U_g2095B (.ZN(g2095B),.A(g143B));
INV_X1 U_g2208B (.ZN(g2208B),.A(g84B));
INV_X1 U_g2579B (.ZN(g2579B),.A(g1969B));
INV_X1 U_I14326B (.ZN(I14326B),.A(g8818B));
INV_X1 U_g6283B (.ZN(g6283B),.A(I9311B));
INV_X1 U_g6920B (.ZN(g6920B),.A(I7817B));
INV_X1 U_g8095B (.ZN(g8095B),.A(g7942B));
INV_X1 U_g6718B (.ZN(g6718B),.A(FE_OFN116_g4807B));
INV_X1 U_g2364B (.ZN(g2364B),.A(g611B));
INV_X1 U_g4194B (.ZN(g4194B),.A(I5399B));
INV_X1 U_g2054B (.ZN(g2054B),.A(g1864B));
INV_X1 U_g6261B (.ZN(g6261B),.A(I9265B));
INV_X1 U_g2725B (.ZN(g2725B),.A(g2018B));
INV_X1 U_g5503B (.ZN(g5503B),.A(FE_OFN204_g3664B));
INV_X1 U_g10465B (.ZN(g10465B),.A(I15986B));
INV_X1 U_g1980B (.ZN(g1980B),.A(g646B));
INV_X1 U_g8164B (.ZN(g8164B),.A(g2216B));
INV_X1 U_g8233B (.ZN(g8233B),.A(g2216B));
INV_X1 U_I6220B (.ZN(I6220B),.A(g883B));
INV_X1 U_I4891B (.ZN(I4891B),.A(g582B));
INV_X1 U_I4859B (.ZN(I4859B),.A(g578B));
INV_X1 U_g4212B (.ZN(g4212B),.A(I5044B));
INV_X1 U_I9479B (.ZN(I9479B),.A(g29B));
INV_X1 U_g2297B (.ZN(g2297B),.A(g865B));
INV_X1 U_g7622B (.ZN(g7622B),.A(g7067B));
INV_X1 U_I13400B (.ZN(I13400B),.A(g8236B));
INV_X1 U_g2338B (.ZN(g2338B),.A(g1909B));
INV_X1 U_g7446B (.ZN(g7446B),.A(FE_OFN86_g2176B));
INV_X1 U_g3475B (.ZN(g3475B),.A(g3056B));
INV_X1 U_g4822B (.ZN(g4822B),.A(g3706B));
INV_X1 U_g10437B (.ZN(g10437B),.A(g10333B));
INV_X1 U_g3039B (.ZN(g3039B),.A(g2310B));
INV_X1 U_I6240B (.ZN(I6240B),.A(g878B));
INV_X1 U_I9810B (.ZN(I9810B),.A(g5576B));
INV_X1 U_g2449B (.ZN(g2449B),.A(g790B));
INV_X1 U_I4783B (.ZN(I4783B),.A(g873B));
INV_X1 U_g2604B (.ZN(g2604B),.A(I5525B));
INV_X1 U_I5399B (.ZN(I5399B),.A(g895B));
INV_X1 U_g6165B (.ZN(g6165B),.A(FE_OFN100_g4421B));
INV_X1 U_I5510B (.ZN(I5510B),.A(g588B));
INV_X1 U_I5245B (.ZN(I5245B),.A(g925B));
INV_X1 U_g9505B (.ZN(g9505B),.A(FE_OFN56_g9052B));
INV_X1 U_g2268B (.ZN(g2268B),.A(g654B));
INV_X1 U_g4192B (.ZN(g4192B),.A(I5388B));
INV_X1 U_g3546B (.ZN(g3546B),.A(FE_OFN352_g109B));
INV_X4 U_g9474B (.ZN(g9474B),.A(g9331B));
INV_X1 U_g5222B (.ZN(g5222B),.A(FE_OFN153_g4640B));
INV_X1 U_g2070B (.ZN(g2070B),.A(g213B));
INV_X1 U_g3906B (.ZN(g3906B),.A(FE_OFN364_g3015B));
INV_X1 U_I4866B (.ZN(I4866B),.A(g579B));
INV_X1 U_g6256B (.ZN(g6256B),.A(g2216B));
INV_X1 U_g4176B (.ZN(g4176B),.A(g1989B));
INV_X1 U_g2331B (.ZN(g2331B),.A(g658B));
INV_X1 U_g2406B (.ZN(g2406B),.A(g1365B));
INV_X1 U_I13332B (.ZN(I13332B),.A(g8206B));
INV_X1 U_g6263B (.ZN(g6263B),.A(I9290B));
INV_X1 U_g11239B (.ZN(g11239B),.A(FE_OFN13_g10702B));
INV_X1 U_g2087B (.ZN(g2087B),.A(g225B));
INV_X1 U_g2801B (.ZN(g2801B),.A(g2117B));
INV_X1 U_g3738B (.ZN(g3738B),.A(g3062B));
INV_X1 U_g7512B (.ZN(g7512B),.A(FE_OFN86_g2176B));
INV_X1 U_g9760B (.ZN(g9760B),.A(FE_OFN33_g9454B));
INV_X1 U_g6257B (.ZN(g6257B),.A(g2169B));
INV_X1 U_g4177B (.ZN(g4177B),.A(g1990B));
INV_X1 U_g4206B (.ZN(g4206B),.A(I5579B));
INV_X1 U_g2045B (.ZN(g2045B),.A(g1811B));
INV_X1 U_g8331B (.ZN(g8331B),.A(I13373B));
INV_X1 U_I9276B (.ZN(I9276B),.A(g83B));
INV_X1 U_g8105B (.ZN(g8105B),.A(g7992B));
INV_X1 U_g2169B (.ZN(g2169B),.A(g42B));
INV_X1 U_I5395B (.ZN(I5395B),.A(g892B));
INV_X1 U_g2369B (.ZN(g2369B),.A(g617B));
INV_X1 U_g2602B (.ZN(g2602B),.A(I5497B));
INV_X1 U_g4199B (.ZN(g4199B),.A(I5418B));
INV_X1 U_g2407B (.ZN(g2407B),.A(g197B));
INV_X1 U_g9451B (.ZN(g9451B),.A(I14642B));
INV_X1 U_g5836B (.ZN(g5836B),.A(FE_OFN273_g85B));
INV_X1 U_g4207B (.ZN(g4207B),.A(I5584B));
INV_X1 U_g11083B (.ZN(g11083B),.A(g10788B));
INV_X1 U_g11348B (.ZN(g11348B),.A(g11276B));
INV_X1 U_I5815B (.ZN(I5815B),.A(g794B));
INV_X1 U_g9508B (.ZN(g9508B),.A(g9271B));
INV_X1 U_g2203B (.ZN(g2203B),.A(g677B));
INV_X1 U_g7686B (.ZN(g7686B),.A(FE_OFN85_g2176B));
INV_X1 U_I5497B (.ZN(I5497B),.A(g587B));
INV_X1 U_I13421B (.ZN(I13421B),.A(g8200B));
INV_X1 U_g4215B (.ZN(g4215B),.A(I5060B));
INV_X1 U_g6863B (.ZN(g6863B),.A(g6740B));
INV_X1 U_g2216B (.ZN(g2216B),.A(g41B));
INV_X1 U_g2028B (.ZN(g2028B),.A(g1703B));
INV_X1 U_g4336B (.ZN(g4336B),.A(g4130B));
INV_X1 U_g2564B (.ZN(g2564B),.A(g1814B));
INV_X1 U_g3705B (.ZN(g3705B),.A(FE_OFN308_I6424B));
INV_X1 U_g4065B (.ZN(g4065B),.A(g2794B));
INV_X1 U_g4887B (.ZN(g4887B),.A(I5057B));
INV_X1 U_g2609B (.ZN(g2609B),.A(I4900B));
INV_X1 U_g4934B (.ZN(g4934B),.A(g4243B));
INV_X1 U_g3814B (.ZN(g3814B),.A(g2355B));
INV_X1 U_g8564B (.ZN(g8564B),.A(I7840B));
INV_X1 U_g2571B (.ZN(g2571B),.A(g1822B));
INV_X1 U_g4195B (.ZN(g4195B),.A(I5406B));
INV_X1 U_g1975B (.ZN(g1975B),.A(g622B));
INV_X1 U_g2774B (.ZN(g2774B),.A(FE_OFN225_g2276B));
INV_X1 U_g3967B (.ZN(g3967B),.A(g3247B));
INV_X1 U_I4935B (.ZN(I4935B),.A(g585B));
INV_X1 U_g2396B (.ZN(g2396B),.A(g1389B));
INV_X1 U_g1984B (.ZN(g1984B),.A(g758B));
INV_X1 U_g11539B (.ZN(g11539B),.A(g11519B));
INV_X1 U_g2018B (.ZN(g2018B),.A(g1336B));
INV_X1 U_g2067B (.ZN(g2067B),.A(g108B));
INV_X1 U_I14323B (.ZN(I14323B),.A(g8817B));
INV_X1 U_I14299B (.ZN(I14299B),.A(g8810B));
INV_X1 U_I6277B (.ZN(I6277B),.A(g1206B));
INV_X1 U_I9237B (.ZN(I9237B),.A(g31B));
INV_X1 U_g2381B (.ZN(g2381B),.A(g1368B));
INV_X1 U_g9432B (.ZN(g9432B),.A(g9313B));
INV_X1 U_g8509B (.ZN(g8509B),.A(g8366B));
INV_X1 U_g7905B (.ZN(g7905B),.A(g7450B));
INV_X1 U_g2421B (.ZN(g2421B),.A(g1374B));
INV_X1 U_g4001B (.ZN(g4001B),.A(g3200B));
INV_X1 U_g11515B (.ZN(g11515B),.A(g11490B));
INV_X1 U_g3485B (.ZN(g3485B),.A(g1104B));
INV_X1 U_g2562B (.ZN(g2562B),.A(g1383B));
INV_X1 U_g6697B (.ZN(g6697B),.A(g4807B));
INV_X1 U_g8700B (.ZN(g8700B),.A(g8574B));
INV_X1 U_g2605B (.ZN(g2605B),.A(I4866B));
INV_X1 U_g11206B (.ZN(g11206B),.A(g10629B));
INV_X1 U_I5427B (.ZN(I5427B),.A(g913B));
INV_X1 U_I9769B (.ZN(I9769B),.A(g5287B));
INV_X1 U_g11107B (.ZN(g11107B),.A(FE_OFN7_g10702B));
INV_X1 U_I11360B (.ZN(I11360B),.A(g6351B));
INV_X1 U_g8562B (.ZN(g8562B),.A(I7825B));
INV_X1 U_g9778B (.ZN(g9778B),.A(FE_OFN63_g9474B));
INV_X1 U_g3765B (.ZN(g3765B),.A(g3120B));
INV_X1 U_g4198B (.ZN(g4198B),.A(I5414B));
INV_X1 U_I14330B (.ZN(I14330B),.A(g8819B));
INV_X1 U_g9526B (.ZN(g9526B),.A(g9256B));
INV_X1 U_I15962B (.ZN(I15962B),.A(g10405B));
INV_X1 U_g3069B (.ZN(g3069B),.A(I6277B));
INV_X1 U_I15500B (.ZN(I15500B),.A(g10019B));
INV_X1 U_I5047B (.ZN(I5047B),.A(g1185B));
INV_X1 U_g2074B (.ZN(g2074B),.A(g1377B));
INV_X1 U_I16507B (.ZN(I16507B),.A(g10712B));
INV_X1 U_g6942B (.ZN(g6942B),.A(I7840B));
INV_X1 U_g4211B (.ZN(g4211B),.A(I5041B));
INV_X1 U_g6432B (.ZN(g6432B),.A(FE_OFN219_g5557B));
INV_X1 U_g7908B (.ZN(g7908B),.A(g7454B));
INV_X1 U_g9764B (.ZN(g9764B),.A(FE_OFN59_g9432B));
INV_X1 U_g3291B (.ZN(g3291B),.A(g2161B));
INV_X1 U_g3207B (.ZN(g3207B),.A(g2439B));
INV_X1 U_g2126B (.ZN(g2126B),.A(g12B));
INV_X1 U_I15514B (.ZN(I15514B),.A(g10007B));
INV_X1 U_I15507B (.ZN(I15507B),.A(g10001B));
INV_X1 U_g1964B (.ZN(g1964B),.A(g114B));
INV_X1 U_g10387B (.ZN(g10387B),.A(g10357B));
INV_X1 U_g11163B (.ZN(g11163B),.A(I16717B));
INV_X1 U_g8688B (.ZN(g8688B),.A(g8507B));
INV_X1 U_g8976B (.ZN(g8976B),.A(I14323B));
INV_X1 U_g2608B (.ZN(g2608B),.A(I4891B));
INV_X1 U_g7450B (.ZN(g7450B),.A(FE_OFN87_g2176B));
INV_X1 U_g4200B (.ZN(g4200B),.A(I5424B));
INV_X1 U_g2023B (.ZN(g2023B),.A(g1357B));
INV_X1 U_g7379B (.ZN(g7379B),.A(g6863B));
INV_X1 U_I13427B (.ZN(I13427B),.A(g8241B));
INV_X1 U_I7752B (.ZN(I7752B),.A(g3407B));
INV_X1 U_g4191B (.ZN(g4191B),.A(I5383B));
INV_X1 U_g1989B (.ZN(g1989B),.A(g770B));
INV_X1 U_g3408B (.ZN(g3408B),.A(g3108B));
INV_X1 U_g2451B (.ZN(g2451B),.A(g248B));
INV_X1 U_g8220B (.ZN(g8220B),.A(FE_OFN199_g7697B));
INV_X1 U_g3943B (.ZN(g3943B),.A(g627B));
INV_X1 U_I14295B (.ZN(I14295B),.A(g8806B));
INV_X1 U_g7981B (.ZN(g7981B),.A(g7624B));
INV_X1 U_g6949B (.ZN(g6949B),.A(I7847B));
INV_X1 U_g8977B (.ZN(g8977B),.A(I14295B));
INV_X1 U_g9082B (.ZN(g9082B),.A(FE_OFN76_g8700B));
INV_X1 U_g4811B (.ZN(g4811B),.A(g3661B));
INV_X1 U_g10379B (.ZN(g10379B),.A(I15861B));
INV_X1 U_g7680B (.ZN(g7680B),.A(FE_OFN87_g2176B));
INV_X1 U_g8327B (.ZN(g8327B),.A(g8164B));
INV_X1 U_I13385B (.ZN(I13385B),.A(g8230B));
INV_X1 U_g7744B (.ZN(g7744B),.A(g1962B));
INV_X1 U_g8146B (.ZN(g8146B),.A(FE_OFN330_g7638B));
INV_X1 U_I5057B (.ZN(I5057B),.A(g1961B));
INV_X1 U_I8503B (.ZN(I8503B),.A(FE_OFN184_I7048B));
INV_X1 U_g2034B (.ZN(g2034B),.A(g1766B));
INV_X1 U_g8103B (.ZN(g8103B),.A(g7994B));
INV_X1 U_g2434B (.ZN(g2434B),.A(g1362B));
INV_X1 U_g3913B (.ZN(g3913B),.A(g3121B));
INV_X1 U_g6702B (.ZN(g6702B),.A(FE_OFN117_g4807B));
INV_X1 U_g4880B (.ZN(g4880B),.A(FE_OFN292_g3015B));
INV_X1 U_g8696B (.ZN(g8696B),.A(g8488B));
INV_X1 U_I14309B (.ZN(I14309B),.A(g8813B));
INV_X1 U_g2347B (.ZN(g2347B),.A(g1945B));
INV_X1 U_g6276B (.ZN(g6276B),.A(I9329B));
INV_X1 U_g4243B (.ZN(g4243B),.A(g3524B));
INV_X1 U_I9259B (.ZN(I9259B),.A(g89B));
INV_X1 U_g7574B (.ZN(g7574B),.A(FE_OFN80_g2175B));
INV_X1 U_g8316B (.ZN(g8316B),.A(I13332B));
INV_X1 U_g8565B (.ZN(g8565B),.A(I7847B));
INV_X1 U_g8347B (.ZN(g8347B),.A(I13421B));
INV_X1 U_g1962B (.ZN(g1962B),.A(g27B));
INV_X1 U_g2601B (.ZN(g2601B),.A(I4859B));
INV_X1 U_g4213B (.ZN(g4213B),.A(I5047B));
INV_X1 U_g6277B (.ZN(g6277B),.A(I9349B));
INV_X1 U_g2060B (.ZN(g2060B),.A(g1380B));
INV_X1 U_g6617B (.ZN(g6617B),.A(g6019B));
INV_X1 U_I13338B (.ZN(I13338B),.A(g8210B));
INV_X1 U_I15861B (.ZN(I15861B),.A(g10339B));
INV_X1 U_I5525B (.ZN(I5525B),.A(g589B));
INV_X1 U_g4456B (.ZN(g4456B),.A(FE_OFN234_g2024B));
INV_X1 U_g2479B (.ZN(g2479B),.A(g26B));
INV_X1 U_I16220B (.ZN(I16220B),.A(g10502B));
INV_X1 U_g9814B (.ZN(g9814B),.A(FE_OFN70_g9490B));
INV_X1 U_g3068B (.ZN(g3068B),.A(g2303B));
INV_X1 U_g9773B (.ZN(g9773B),.A(g9474B));
INV_X1 U_g5200B (.ZN(g5200B),.A(g4567B));
INV_X1 U_g4457B (.ZN(g4457B),.A(FE_OFN137_g3829B));
INV_X1 U_g4193B (.ZN(g4193B),.A(I5395B));
INV_X1 U_g10461B (.ZN(g10461B),.A(I15974B));
INV_X1 U_I5020B (.ZN(I5020B),.A(g1176B));
INV_X1 U_g1969B (.ZN(g1969B),.A(g456B));
INV_X1 U_I9293B (.ZN(I9293B),.A(g92B));
INV_X1 U_I9329B (.ZN(I9329B),.A(g94B));
INV_X1 U_g7903B (.ZN(g7903B),.A(g7446B));
INV_X1 U_I9221B (.ZN(I9221B),.A(g30B));
INV_X1 U_g4525B (.ZN(g4525B),.A(FE_OFN229_g3880B));
INV_X1 U_g2475B (.ZN(g2475B),.A(g192B));
INV_X1 U_g1988B (.ZN(g1988B),.A(g766B));
INV_X1 U_g11203B (.ZN(g11203B),.A(FE_OFN20_g10702B));
INV_X1 U_g4158B (.ZN(g4158B),.A(g3304B));
INV_X1 U_g6557B (.ZN(g6557B),.A(FE_OFN217_g5013B));
INV_X1 U_g2603B (.ZN(g2603B),.A(I5510B));
INV_X1 U_I5410B (.ZN(I5410B),.A(g901B));
INV_X1 U_g10459B (.ZN(g10459B),.A(I15968B));
INV_X1 U_I9349B (.ZN(I9349B),.A(g95B));
INV_X1 U_g6955B (.ZN(g6955B),.A(I7852B));
INV_X1 U_I15290B (.ZN(I15290B),.A(g9974B));
INV_X1 U_g6254B (.ZN(g6254B),.A(I9221B));
INV_X1 U_g4174B (.ZN(g4174B),.A(g1987B));
INV_X1 U_g10444B (.ZN(g10444B),.A(g10325B));
INV_X1 U_I14642B (.ZN(I14642B),.A(g9088B));
INV_X1 U_g4180B (.ZN(g4180B),.A(g1993B));
INV_X1 U_g7917B (.ZN(g7917B),.A(g7497B));
INV_X1 U_g2986B (.ZN(g2986B),.A(I6220B));
INV_X1 U_g9473B (.ZN(g9473B),.A(g9082B));
INV_X1 U_g1965B (.ZN(g1965B),.A(g119B));
INV_X1 U_g11547B (.ZN(g11547B),.A(FE_OFN27_g11519B));
INV_X1 U_g2503B (.ZN(g2503B),.A(g1872B));
INV_X1 U_I9352B (.ZN(I9352B),.A(g28B));
INV_X1 U_I9717B (.ZN(I9717B),.A(FE_OFN97_I8869B));
INV_X1 U_g2224B (.ZN(g2224B),.A(g695B));
INV_X1 U_g7454B (.ZN(g7454B),.A(g2176B));
INV_X1 U_g4204B (.ZN(g4204B),.A(I5445B));
INV_X1 U_g8561B (.ZN(g8561B),.A(I7817B));
INV_X1 U_g8986B (.ZN(g8986B),.A(I14330B));
INV_X1 U_I15956B (.ZN(I15956B),.A(g10402B));
INV_X1 U_I15980B (.ZN(I15980B),.A(g10414B));
AND2_X1 U_g11103B (.ZN(g11103B),.A2(g10937B),.A1(g2250B));
AND2_X1 U_g9900B (.ZN(g9900B),.A2(g8327B),.A1(g9088B));
AND2_X1 U_g11095B (.ZN(g11095B),.A2(FE_OFN4_g10950B),.A1(g845B));
AND2_X2 U_g3880B (.ZN(g3880B),.A2(g2023B),.A1(FE_OFN235_g2024B));
AND2_X1 U_g4973B (.ZN(g4973B),.A2(g4467B),.A1(g1645B));
AND2_X1 U_g7389B (.ZN(g7389B),.A2(FE_OFN226_g3880B),.A1(g5852B));
AND2_X1 U_g7888B (.ZN(g7888B),.A2(FE_OFN334_g7045B),.A1(g7465B));
AND2_X1 U_g4969B (.ZN(g4969B),.A2(g4457B),.A1(g1642B));
AND2_X1 U_g8224B (.ZN(g8224B),.A2(g7949B),.A1(g1882B));
AND2_X1 U_g2892B (.ZN(g2892B),.A2(g1976B),.A1(g1980B));
AND2_X1 U_g5686B (.ZN(g5686B),.A2(FE_OFN365_g5361B),.A1(g158B));
AND2_X1 U_g10308B (.ZN(g10308B),.A2(g9082B),.A1(g10013B));
AND2_X1 U_g4123B (.ZN(g4123B),.A2(g2424B),.A1(g1781B));
AND2_X1 U_g8120B (.ZN(g8120B),.A2(g7949B),.A1(g1909B));
AND2_X1 U_g6788B (.ZN(g6788B),.A2(FE_OFN320_g5361B),.A1(g287B));
AND2_X1 U_g5598B (.ZN(g5598B),.A2(g4824B),.A1(g778B));
AND2_X1 U_g9694B (.ZN(g9694B),.A2(FE_OFN59_g9432B),.A1(g278B));
AND2_X1 U_g10495B (.ZN(g10495B),.A2(FE_OFN234_g2024B),.A1(g10431B));
AND2_X1 U_g2945B (.ZN(g2945B),.A2(g1684B),.A1(FE_OFN241_g1690B));
AND2_X1 U_g11190B (.ZN(g11190B),.A2(g10927B),.A1(g4752B));
AND2_X1 U_g8789B (.ZN(g8789B),.A2(FE_OFN331_g8696B),.A1(g8639B));
AND2_X1 U_g9852B (.ZN(g9852B),.A2(g9563B),.A1(g9728B));
AND2_X1 U_g5625B (.ZN(g5625B),.A2(g5627B),.A1(g1053B));
AND2_X1 U_g4875B (.ZN(g4875B),.A2(g4673B),.A1(g995B));
AND2_X1 U_g9701B (.ZN(g9701B),.A2(g9474B),.A1(g1574B));
AND2_X1 U_g7138B (.ZN(g7138B),.A2(g6718B),.A1(g5201B));
AND2_X1 U_g10752B (.ZN(g10752B),.A2(FE_OFN103_g3586B),.A1(g10599B));
AND2_X1 U_g11211B (.ZN(g11211B),.A2(g5503B),.A1(g11058B));
AND2_X1 U_g11024B (.ZN(g11024B),.A2(g10702B),.A1(g435B));
AND2_X1 U_g8547B (.ZN(g8547B),.A2(FE_OFN211_g7246B),.A1(g8307B));
AND2_X1 U_g10669B (.ZN(g10669B),.A2(g9473B),.A1(g10408B));
AND2_X1 U_g7707B (.ZN(g7707B),.A2(FE_OFN191_g6488B),.A1(g691B));
AND2_X1 U_g4884B (.ZN(g4884B),.A2(g1845B),.A1(g3813B));
AND2_X1 U_g4839B (.ZN(g4839B),.A2(g2355B),.A1(g225B));
AND2_X1 U_g9870B (.ZN(g9870B),.A2(g9802B),.A1(g1561B));
AND2_X1 U_g6640B (.ZN(g6640B),.A2(g5808B),.A1(g86B));
AND2_X1 U_g9650B (.ZN(g9650B),.A2(FE_OFN40_g9240B),.A1(g986B));
AND2_X1 U_g5687B (.ZN(g5687B),.A2(FE_OFN365_g5361B),.A1(g139B));
AND2_X1 U_g7957B (.ZN(g7957B),.A2(g7527B),.A1(g79B));
AND2_X1 U_g3512B (.ZN(g3512B),.A2(g1845B),.A1(g2050B));
AND2_X1 U_g8244B (.ZN(g8244B),.A2(FE_OFN310_g4336B),.A1(g7054B));
AND2_X1 U_g7449B (.ZN(g7449B),.A2(FE_OFN221_g3440B),.A1(g6548B));
AND2_X1 U_g4235B (.ZN(g4235B),.A2(FE_OFN347_g3914B),.A1(g1011B));
AND2_X1 U_g4343B (.ZN(g4343B),.A2(FE_OFN287_g3586B),.A1(g345B));
AND2_X1 U_g11296B (.ZN(g11296B),.A2(g11239B),.A1(g4561B));
AND2_X1 U_g9594B (.ZN(g9594B),.A2(g9292B),.A1(g1B));
AND2_X1 U_g6829B (.ZN(g6829B),.A2(FE_OFN179_g5354B),.A1(g213B));
AND2_X1 U_g4334B (.ZN(g4334B),.A2(FE_OFN351_g3913B),.A1(g1160B));
AND2_X1 U_g9943B (.ZN(g9943B),.A2(FE_OFN67_g9367B),.A1(g9923B));
AND2_X1 U_g5525B (.ZN(g5525B),.A2(g4292B),.A1(g1721B));
AND2_X1 U_g4548B (.ZN(g4548B),.A2(g4002B),.A1(g440B));
AND3_X1 U_g8876B (.ZN(g8876B),.A3(FE_OFN73_g8858B),.A2(FE_OFN93_g2216B),.A1(g8105B));
AND2_X1 U_g6733B (.ZN(g6733B),.A2(FE_OFN322_g4449B),.A1(g4488B));
AND2_X1 U_g4804B (.ZN(g4804B),.A2(g4010B),.A1(g476B));
AND2_X1 U_g10705B (.ZN(g10705B),.A2(FE_OFN131_g3015B),.A1(g10564B));
AND2_X1 U_g9934B (.ZN(g9934B),.A2(g9624B),.A1(g9913B));
AND2_X1 U_g6225B (.ZN(g6225B),.A2(g5613B),.A1(g566B));
AND2_X1 U_g6324B (.ZN(g6324B),.A2(FE_OFN116_g4807B),.A1(g1240B));
AND2_X1 U_g10686B (.ZN(g10686B),.A2(FE_OFN136_g3863B),.A1(g10385B));
AND2_X1 U_g6540B (.ZN(g6540B),.A2(g6081B),.A1(g1223B));
AND2_X1 U_g8663B (.ZN(g8663B),.A2(FE_OFN292_g3015B),.A1(g8270B));
AND2_X1 U_g11581B (.ZN(g11581B),.A2(g11539B),.A1(g1308B));
AND2_X1 U_g6206B (.ZN(g6206B),.A2(g5613B),.A1(g560B));
AND2_X1 U_g4518B (.ZN(g4518B),.A2(g4002B),.A1(g452B));
AND2_X1 U_g3989B (.ZN(g3989B),.A2(FE_OFN359_g18B),.A1(g248B));
AND2_X1 U_g7730B (.ZN(g7730B),.A2(g2347B),.A1(g7260B));
AND2_X1 U_g5174B (.ZN(g5174B),.A2(FE_OFN303_g4678B),.A1(g1235B));
AND2_X1 U_g7504B (.ZN(g7504B),.A2(g67B),.A1(FE_OFN86_g2176B));
AND2_X1 U_g7185B (.ZN(g7185B),.A2(FE_OFN213_g6003B),.A1(g1887B));
AND2_X1 U_g2563B (.ZN(g2563B),.A2(I5690B),.A1(I5689B));
AND2_X1 U_g7881B (.ZN(g7881B),.A2(FE_OFN366_g3521B),.A1(g5295B));
AND2_X1 U_g11070B (.ZN(g11070B),.A2(g10788B),.A1(g2008B));
AND2_X1 U_g9859B (.ZN(g9859B),.A2(g9579B),.A1(g9736B));
AND3_X1 U_g8877B (.ZN(g8877B),.A3(FE_OFN73_g8858B),.A2(FE_OFN92_g2216B),.A1(g8103B));
AND2_X1 U_g11590B (.ZN(g11590B),.A2(g11561B),.A1(g2274B));
AND2_X1 U_g6199B (.ZN(g6199B),.A2(FE_OFN289_g4679B),.A1(g557B));
AND2_X1 U_g9266B (.ZN(g9266B),.A2(FE_OFN325_g18B),.A1(g8932B));
AND2_X1 U_g5545B (.ZN(g5545B),.A2(g4292B),.A1(g1730B));
AND2_X1 U_g5180B (.ZN(g5180B),.A2(g810B),.A1(g814B));
AND2_X1 U_g5591B (.ZN(g5591B),.A2(FE_OFN367_g3521B),.A1(g1615B));
AND2_X1 U_g8556B (.ZN(g8556B),.A2(FE_OFN189_g7638B),.A1(g8412B));
AND2_X1 U_g11094B (.ZN(g11094B),.A2(g10883B),.A1(g374B));
AND2_X1 U_g5853B (.ZN(g5853B),.A2(g1927B),.A1(g5044B));
AND2_X1 U_g6245B (.ZN(g6245B),.A2(FE_OFN289_g4679B),.A1(g575B));
AND2_X1 U_g4360B (.ZN(g4360B),.A2(g3523B),.A1(g1861B));
AND3_X1 U_g8930B (.ZN(g8930B),.A3(g8828B),.A2(FE_OFN95_g2216B),.A1(g8100B));
AND2_X1 U_g5507B (.ZN(g5507B),.A2(FE_OFN357_g3521B),.A1(g563B));
AND2_X1 U_g11150B (.ZN(g11150B),.A2(g10788B),.A1(g3087B));
AND2_X1 U_g8464B (.ZN(g8464B),.A2(FE_OFN210_g7246B),.A1(g8302B));
AND2_X1 U_g9692B (.ZN(g9692B),.A2(FE_OFN59_g9432B),.A1(g272B));
AND2_X1 U_g4996B (.ZN(g4996B),.A2(FE_OFN146_g4682B),.A1(g1428B));
AND2_X1 U_g7131B (.ZN(g7131B),.A2(g6702B),.A1(g5174B));
AND2_X1 U_g11019B (.ZN(g11019B),.A2(FE_OFN7_g10702B),.A1(g421B));
AND2_X1 U_g9960B (.ZN(g9960B),.A2(FE_OFN280_g9536B),.A1(g9951B));
AND2_X1 U_g11196B (.ZN(g11196B),.A2(FE_OFN15_g10702B),.A1(g4770B));
AND2_X1 U_g11018B (.ZN(g11018B),.A2(FE_OFN7_g10702B),.A1(g6485B));
AND2_X1 U_g6819B (.ZN(g6819B),.A2(FE_OFN179_g5354B),.A1(g243B));
AND2_X1 U_g10595B (.ZN(g10595B),.A2(FE_OFN369_g4525B),.A1(g10550B));
AND2_X1 U_g10494B (.ZN(g10494B),.A2(g2024B),.A1(g10433B));
AND2_X1 U_g10623B (.ZN(g10623B),.A2(FE_OFN370_g4525B),.A1(g10544B));
AND2_X1 U_g4878B (.ZN(g4878B),.A2(g3523B),.A1(g1868B));
AND2_X1 U_g5204B (.ZN(g5204B),.A2(g2126B),.A1(g4838B));
AND2_X1 U_g8844B (.ZN(g8844B),.A2(g8709B),.A1(g8609B));
AND2_X1 U_g6701B (.ZN(g6701B),.A2(g4381B),.A1(g6185B));
AND2_X1 U_g10782B (.ZN(g10782B),.A2(g4467B),.A1(g10725B));
AND2_X1 U_g5100B (.ZN(g5100B),.A2(g4608B),.A1(g1791B));
AND2_X1 U_g4882B (.ZN(g4882B),.A2(FE_OFN293_g3015B),.A1(g1089B));
AND2_X1 U_g8731B (.ZN(g8731B),.A2(g7918B),.A1(g8236B));
AND2_X1 U_g6215B (.ZN(g6215B),.A2(g5128B),.A1(g1504B));
AND2_X1 U_g6886B (.ZN(g6886B),.A2(FE_OFN213_g6003B),.A1(g1932B));
AND2_X4 U_g3586B (.ZN(g3586B),.A2(I6260B),.A1(g1703B));
AND2_X1 U_g8557B (.ZN(g8557B),.A2(g7638B),.A1(g8415B));
AND3_X1 U_g8966B (.ZN(g8966B),.A3(g8849B),.A2(FE_OFN93_g2216B),.A1(g8081B));
AND2_X1 U_g8071B (.ZN(g8071B),.A2(FE_OFN199_g7697B),.A1(g691B));
AND2_X1 U_g11597B (.ZN(g11597B),.A2(FE_OFN99_g4421B),.A1(g11549B));
AND2_X1 U_g9828B (.ZN(g9828B),.A2(g9785B),.A1(g9722B));
AND2_X1 U_g2918B (.ZN(g2918B),.A2(g1672B),.A1(FE_OFN241_g1690B));
AND2_X1 U_g9830B (.ZN(g9830B),.A2(FE_OFN34_g9785B),.A1(g9725B));
AND3_X1 U_g8955B (.ZN(g8955B),.A3(g8828B),.A2(FE_OFN95_g2216B),.A1(g8110B));
AND2_X1 U_g9592B (.ZN(g9592B),.A2(g9292B),.A1(g4B));
AND2_X1 U_g5123B (.ZN(g5123B),.A2(g3906B),.A1(g1618B));
AND2_X1 U_g7059B (.ZN(g7059B),.A2(g6354B),.A1(g6078B));
AND2_X1 U_g8254B (.ZN(g8254B),.A2(g7907B),.A1(g936B));
AND2_X1 U_g7459B (.ZN(g7459B),.A2(g55B),.A1(FE_OFN86_g2176B));
AND2_X1 U_g11102B (.ZN(g11102B),.A2(FE_OFN3_g10950B),.A1(g861B));
AND2_X1 U_g7718B (.ZN(g7718B),.A2(FE_OFN191_g6488B),.A1(g709B));
AND2_X1 U_g7535B (.ZN(g7535B),.A2(g49B),.A1(FE_OFN86_g2176B));
AND2_X1 U_g9703B (.ZN(g9703B),.A2(g9474B),.A1(g1577B));
AND2_X1 U_g5528B (.ZN(g5528B),.A2(FE_OFN357_g3521B),.A1(g569B));
AND2_X1 U_g9932B (.ZN(g9932B),.A2(g9624B),.A1(g9911B));
AND2_X1 U_g5530B (.ZN(g5530B),.A2(FE_OFN290_g4880B),.A1(g1636B));
AND2_X1 U_g3506B (.ZN(g3506B),.A2(g2760B),.A1(g986B));
AND2_X1 U_g8769B (.ZN(g8769B),.A2(FE_OFN304_g5151B),.A1(g8629B));
AND2_X1 U_g6887B (.ZN(g6887B),.A2(g6557B),.A1(g6187B));
AND2_X1 U_g6228B (.ZN(g6228B),.A2(g713B),.A1(g5605B));
AND2_X1 U_g6322B (.ZN(g6322B),.A2(FE_OFN116_g4807B),.A1(g1275B));
AND2_X1 U_g3111B (.ZN(g3111B),.A2(I6338B),.A1(I6337B));
AND3_X1 U_g8967B (.ZN(g8967B),.A3(g8849B),.A2(FE_OFN281_g2216B),.A1(g8085B));
AND2_X1 U_g5010B (.ZN(g5010B),.A2(FE_OFN153_g4640B),.A1(g1458B));
AND2_X1 U_g3275B (.ZN(g3275B),.A2(FE_OFN266_g18B),.A1(g115B));
AND2_X1 U_g10809B (.ZN(g10809B),.A2(g10702B),.A1(g4811B));
AND2_X1 U_g2895B (.ZN(g2895B),.A2(g1678B),.A1(FE_OFN336_g1690B));
AND2_X1 U_g7721B (.ZN(g7721B),.A2(g6488B),.A1(g736B));
AND2_X1 U_g9866B (.ZN(g9866B),.A2(g9802B),.A1(g1549B));
AND2_X1 U_g9716B (.ZN(g9716B),.A2(FE_OFN70_g9490B),.A1(g1534B));
AND2_X1 U_g10808B (.ZN(g10808B),.A2(FE_OFN137_g3829B),.A1(g10744B));
AND2_X1 U_g3374B (.ZN(g3374B),.A2(g3047B),.A1(g1231B));
AND2_X1 U_g4492B (.ZN(g4492B),.A2(g3685B),.A1(FE_OFN253_g1786B));
AND2_X1 U_g8822B (.ZN(g8822B),.A2(FE_OFN328_g8709B),.A1(g8614B));
AND2_X1 U_g10560B (.ZN(g10560B),.A2(FE_OFN369_g4525B),.A1(g10369B));
AND3_X1 U_g11456B (.ZN(g11456B),.A3(g11348B),.A2(g2801B),.A1(g3765B));
AND2_X1 U_g9848B (.ZN(g9848B),.A2(g9579B),.A1(g9724B));
AND2_X1 U_g4714B (.ZN(g4714B),.A2(g3943B),.A1(g646B));
AND2_X1 U_g6550B (.ZN(g6550B),.A2(g6081B),.A1(g1231B));
AND2_X1 U_g5172B (.ZN(g5172B),.A2(g818B),.A1(g822B));
AND2_X1 U_g10642B (.ZN(g10642B),.A2(g3829B),.A1(g10385B));
AND2_X1 U_g3284B (.ZN(g3284B),.A2(g677B),.A1(g2531B));
AND2_X1 U_g9699B (.ZN(g9699B),.A2(FE_OFN59_g9432B),.A1(g284B));
AND2_X1 U_g9855B (.ZN(g9855B),.A2(g9764B),.A1(g302B));
AND2_X1 U_g5618B (.ZN(g5618B),.A2(FE_OFN367_g3521B),.A1(g1630B));
AND2_X1 U_g6891B (.ZN(g6891B),.A2(g6003B),.A1(g1950B));
AND2_X1 U_g7940B (.ZN(g7940B),.A2(FE_OFN292_g3015B),.A1(g5319B));
AND2_X1 U_g11085B (.ZN(g11085B),.A2(g10927B),.A1(g312B));
AND2_X1 U_g4736B (.ZN(g4736B),.A2(FE_OFN300_g4002B),.A1(g396B));
AND2_X1 U_g4968B (.ZN(g4968B),.A2(FE_OFN146_g4682B),.A1(g1432B));
AND2_X1 U_g8837B (.ZN(g8837B),.A2(FE_OFN331_g8696B),.A1(g8646B));
AND2_X1 U_g9644B (.ZN(g9644B),.A2(FE_OFN45_g9125B),.A1(g1182B));
AND2_X1 U_g5804B (.ZN(g5804B),.A2(g5261B),.A1(g1546B));
AND2_X1 U_g8462B (.ZN(g8462B),.A2(FE_OFN211_g7246B),.A1(g8300B));
AND4_X1 U_I6330B (.ZN(I6330B),.A4(g2570B),.A3(g2562B),.A2(g2556B),.A1(g2549B));
AND2_X1 U_g11156B (.ZN(g11156B),.A2(FE_OFN278_g10927B),.A1(g333B));
AND2_X1 U_g6342B (.ZN(g6342B),.A2(FE_OFN319_g5361B),.A1(g293B));
AND2_X1 U_g9867B (.ZN(g9867B),.A2(g9802B),.A1(g1552B));
AND2_X1 U_g9717B (.ZN(g9717B),.A2(FE_OFN70_g9490B),.A1(g1537B));
AND2_X1 U_g4871B (.ZN(g4871B),.A2(g3523B),.A1(g1864B));
AND2_X1 U_g10454B (.ZN(g10454B),.A2(FE_OFN235_g2024B),.A1(g10435B));
AND2_X1 U_g4722B (.ZN(g4722B),.A2(FE_OFN300_g4002B),.A1(g426B));
AND2_X1 U_g7741B (.ZN(g7741B),.A2(g3880B),.A1(g5824B));
AND2_X1 U_g4500B (.ZN(g4500B),.A2(FE_OFN291_g4880B),.A1(g1357B));
AND2_X1 U_g9386B (.ZN(g9386B),.A2(FE_OFN47_g9151B),.A1(g1327B));
AND2_X1 U_g8842B (.ZN(g8842B),.A2(FE_OFN328_g8709B),.A1(g8607B));
AND2_X1 U_g9599B (.ZN(g9599B),.A2(FE_OFN71_g9292B),.A1(g8B));
AND2_X4 U_g9274B (.ZN(g9274B),.A2(FE_OFN275_g48B),.A1(g8974B));
AND2_X1 U_g5518B (.ZN(g5518B),.A2(FE_OFN357_g3521B),.A1(g566B));
AND2_X1 U_g9614B (.ZN(g9614B),.A2(FE_OFN51_g9111B),.A1(g1197B));
AND2_X1 U_g4838B (.ZN(g4838B),.A2(g4122B),.A1(g3275B));
AND2_X4 U_g9125B (.ZN(g9125B),.A2(FE_OFN276_g48B),.A1(g8966B));
AND2_X1 U_g7217B (.ZN(g7217B),.A2(g6432B),.A1(g4610B));
AND2_X1 U_g11557B (.ZN(g11557B),.A2(g11519B),.A1(g1791B));
AND2_X1 U_g2911B (.ZN(g2911B),.A2(g1675B),.A1(FE_OFN336_g1690B));
AND2_X1 U_g11210B (.ZN(g11210B),.A2(FE_OFN204_g3664B),.A1(g10886B));
AND2_X1 U_g7466B (.ZN(g7466B),.A2(g58B),.A1(g2176B));
AND2_X1 U_g9939B (.ZN(g9939B),.A2(FE_OFN67_g9367B),.A1(g9918B));
AND2_X1 U_g11279B (.ZN(g11279B),.A2(g11203B),.A1(g4784B));
AND3_X1 U_g10518B (.ZN(g10518B),.A3(I16145B),.A2(g10440B),.A1(g10513B));
AND2_X1 U_g4477B (.ZN(g4477B),.A2(g3913B),.A1(g1129B));
AND2_X1 U_g7055B (.ZN(g7055B),.A2(g6586B),.A1(g5004B));
AND2_X1 U_g5264B (.ZN(g5264B),.A2(g4776B),.A1(g1095B));
AND2_X1 U_g6329B (.ZN(g6329B),.A2(FE_OFN115_g4807B),.A1(g1265B));
AND2_X1 U_g6828B (.ZN(g6828B),.A2(FE_OFN179_g5354B),.A1(g1377B));
AND2_X1 U_g8176B (.ZN(g8176B),.A2(FE_OFN89_I11360B),.A1(g40B));
AND2_X1 U_g6830B (.ZN(g6830B),.A2(FE_OFN179_g5354B),.A1(g1380B));
AND2_X1 U_g8005B (.ZN(g8005B),.A2(FE_OFN334_g7045B),.A1(g7510B));
AND2_X1 U_g4099B (.ZN(g4099B),.A2(g3281B),.A1(g770B));
AND2_X1 U_g11601B (.ZN(g11601B),.A2(g11575B),.A1(g1351B));
AND2_X1 U_g11187B (.ZN(g11187B),.A2(FE_OFN10_g10702B),.A1(g4727B));
AND2_X1 U_g6746B (.ZN(g6746B),.A2(FE_OFN218_g5557B),.A1(g6228B));
AND2_X1 U_g6221B (.ZN(g6221B),.A2(g5598B),.A1(g782B));
AND2_X1 U_g8765B (.ZN(g8765B),.A2(FE_OFN304_g5151B),.A1(g8630B));
AND2_X1 U_g9622B (.ZN(g9622B),.A2(FE_OFN51_g9111B),.A1(g1200B));
AND2_X1 U_g11143B (.ZN(g11143B),.A2(g4567B),.A1(g10923B));
AND2_X1 U_g9904B (.ZN(g9904B),.A2(g9676B),.A1(g9886B));
AND2_X1 U_g8733B (.ZN(g8733B),.A2(g7920B),.A1(g8241B));
AND3_X1 U_g8974B (.ZN(g8974B),.A3(FE_OFN73_g8858B),.A2(FE_OFN93_g2216B),.A1(g8094B));
AND2_X1 U_g6624B (.ZN(g6624B),.A2(FE_OFN282_g6165B),.A1(g348B));
AND2_X1 U_g11169B (.ZN(g11169B),.A2(FE_OFN8_g10702B),.A1(g530B));
AND2_X1 U_g8073B (.ZN(g8073B),.A2(FE_OFN199_g7697B),.A1(g709B));
AND2_X1 U_g9841B (.ZN(g9841B),.A2(g9512B),.A1(g9706B));
AND2_X1 U_g5882B (.ZN(g5882B),.A2(FE_OFN141_g3829B),.A1(g5592B));
AND2_X1 U_g8796B (.ZN(g8796B),.A2(FE_OFN331_g8696B),.A1(g8645B));
AND2_X1 U_g11168B (.ZN(g11168B),.A2(FE_OFN7_g10702B),.A1(g534B));
AND2_X1 U_g4269B (.ZN(g4269B),.A2(FE_OFN347_g3914B),.A1(g1015B));
AND2_X1 U_g5271B (.ZN(g5271B),.A2(FE_OFN335_g4737B),.A1(g727B));
AND2_X1 U_g10348B (.ZN(g10348B),.A2(g3705B),.A1(I15500B));
AND2_X1 U_g5611B (.ZN(g5611B),.A2(g4880B),.A1(g1047B));
AND2_X1 U_g8069B (.ZN(g8069B),.A2(FE_OFN198_g7697B),.A1(g673B));
AND2_X1 U_g9695B (.ZN(g9695B),.A2(g9474B),.A1(g1567B));
AND2_X1 U_g10304B (.ZN(g10304B),.A2(g9291B),.A1(g10001B));
AND2_X1 U_g8469B (.ZN(g8469B),.A2(FE_OFN211_g7246B),.A1(g8305B));
AND2_X1 U_g4712B (.ZN(g4712B),.A2(FE_OFN297_g3015B),.A1(g1071B));
AND2_X1 U_g6576B (.ZN(g6576B),.A2(g5503B),.A1(g5762B));
AND2_X1 U_g10622B (.ZN(g10622B),.A2(FE_OFN369_g4525B),.A1(g10496B));
AND2_X1 U_g11015B (.ZN(g11015B),.A2(FE_OFN18_g10702B),.A1(g5217B));
AND2_X1 U_g5674B (.ZN(g5674B),.A2(FE_OFN365_g5361B),.A1(g148B));
AND2_X1 U_g9359B (.ZN(g9359B),.A2(FE_OFN52_g9173B),.A1(g1308B));
AND2_X2 U_g9223B (.ZN(g9223B),.A2(g8960B),.A1(FE_OFN277_g48B));
AND2_X1 U_g11556B (.ZN(g11556B),.A2(g11519B),.A1(g1786B));
AND2_X1 U_g9858B (.ZN(g9858B),.A2(g9778B),.A1(g1595B));
AND2_X1 U_g5541B (.ZN(g5541B),.A2(g3521B),.A1(g575B));
AND2_X1 U_g4534B (.ZN(g4534B),.A2(FE_OFN344_g3586B),.A1(g363B));
AND2_X1 U_g6198B (.ZN(g6198B),.A2(g5128B),.A1(g1499B));
AND2_X1 U_g6747B (.ZN(g6747B),.A2(g5897B),.A1(g2214B));
AND2_X1 U_g6699B (.ZN(g6699B),.A2(FE_OFN111_g3914B),.A1(g6177B));
AND2_X1 U_g6855B (.ZN(g6855B),.A2(g6392B),.A1(g1964B));
AND2_X1 U_g3804B (.ZN(g3804B),.A2(g2203B),.A1(g3098B));
AND2_X1 U_g5680B (.ZN(g5680B),.A2(FE_OFN164_g5361B),.A1(g153B));
AND2_X1 U_g9642B (.ZN(g9642B),.A2(FE_OFN40_g9240B),.A1(g981B));
AND2_X1 U_g5744B (.ZN(g5744B),.A2(FE_OFN321_g5261B),.A1(g1528B));
AND2_X1 U_g10333B (.ZN(g10333B),.A2(FE_OFN267_g109B),.A1(I15500B));
AND2_X1 U_g8399B (.ZN(g8399B),.A2(g8220B),.A1(g5266B));
AND2_X1 U_g9447B (.ZN(g9447B),.A2(FE_OFN49_g9030B),.A1(g1762B));
AND2_X1 U_g4903B (.ZN(g4903B),.A2(g4243B),.A1(g1849B));
AND2_X1 U_g11178B (.ZN(g11178B),.A2(FE_OFN13_g10702B),.A1(g516B));
AND2_X1 U_g8510B (.ZN(g8510B),.A2(FE_OFN330_g7638B),.A1(g8414B));
AND2_X1 U_g8245B (.ZN(g8245B),.A2(FE_OFN322_g4449B),.A1(g7062B));
AND2_X1 U_g6319B (.ZN(g6319B),.A2(FE_OFN118_g4807B),.A1(g1296B));
AND2_X1 U_g11186B (.ZN(g11186B),.A2(FE_OFN10_g10702B),.A1(g4722B));
AND2_X1 U_g2951B (.ZN(g2951B),.A2(g1681B),.A1(FE_OFN241_g1690B));
AND2_X1 U_g6352B (.ZN(g6352B),.A2(FE_OFN319_g5361B),.A1(g278B));
AND2_X1 U_g9595B (.ZN(g9595B),.A2(FE_OFN42_g9205B),.A1(g901B));
AND2_X1 U_g4831B (.ZN(g4831B),.A2(g4109B),.A1(g810B));
AND2_X1 U_g5492B (.ZN(g5492B),.A2(g4263B),.A1(g1654B));
AND2_X1 U_g9272B (.ZN(g9272B),.A2(FE_OFN266_g18B),.A1(g8934B));
AND2_X1 U_g10312B (.ZN(g10312B),.A2(g9082B),.A1(g10019B));
AND2_X1 U_g6186B (.ZN(g6186B),.A2(FE_OFN291_g4880B),.A1(g546B));
AND2_X1 U_g9612B (.ZN(g9612B),.A2(FE_OFN40_g9240B),.A1(g2652B));
AND2_X1 U_g9417B (.ZN(g9417B),.A2(FE_OFN56_g9052B),.A1(g1738B));
AND2_X1 U_g9935B (.ZN(g9935B),.A2(FE_OFN60_g9624B),.A1(g9914B));
AND2_X1 U_g10745B (.ZN(g10745B),.A2(FE_OFN102_g3586B),.A1(g10658B));
AND2_X1 U_g11216B (.ZN(g11216B),.A2(FE_OFN279_g11157B),.A1(g956B));
AND2_X1 U_g9328B (.ZN(g9328B),.A2(FE_OFN275_g48B),.A1(g8971B));
AND2_X1 U_g11587B (.ZN(g11587B),.A2(g11539B),.A1(g1327B));
AND2_X1 U_g6821B (.ZN(g6821B),.A2(FE_OFN178_g5354B),.A1(g237B));
AND2_X1 U_g6325B (.ZN(g6325B),.A2(FE_OFN116_g4807B),.A1(g1245B));
AND2_X1 U_g4560B (.ZN(g4560B),.A2(g4002B),.A1(g431B));
AND2_X1 U_g7368B (.ZN(g7368B),.A2(g3880B),.A1(g5842B));
AND2_X1 U_g6083B (.ZN(g6083B),.A2(g4273B),.A1(g552B));
AND2_X1 U_g6544B (.ZN(g6544B),.A2(g6081B),.A1(g1227B));
AND2_X1 U_g5476B (.ZN(g5476B),.A2(g4673B),.A1(g1615B));
AND2_X1 U_g7743B (.ZN(g7743B),.A2(FE_OFN226_g3880B),.A1(g5838B));
AND2_X1 U_g4869B (.ZN(g4869B),.A2(FE_OFN132_g3015B),.A1(g1083B));
AND2_X1 U_g5722B (.ZN(g5722B),.A2(FE_OFN315_g5117B),.A1(g1598B));
AND2_X1 U_g6790B (.ZN(g6790B),.A2(FE_OFN346_g4381B),.A1(g5813B));
AND2_X1 U_g8408B (.ZN(g8408B),.A2(g8146B),.A1(g704B));
AND2_X1 U_g10761B (.ZN(g10761B),.A2(g10558B),.A1(g10559B));
AND2_X1 U_g7734B (.ZN(g7734B),.A2(FE_OFN226_g3880B),.A1(g5810B));
AND2_X1 U_g8136B (.ZN(g8136B),.A2(g7045B),.A1(g7926B));
AND2_X1 U_g6187B (.ZN(g6187B),.A2(g2340B),.A1(g5569B));
AND2_X1 U_g4752B (.ZN(g4752B),.A2(FE_OFN300_g4002B),.A1(g401B));
AND2_X1 U_g9902B (.ZN(g9902B),.A2(FE_OFN69_g9392B),.A1(g9720B));
AND2_X1 U_g8768B (.ZN(g8768B),.A2(FE_OFN304_g5151B),.A1(g8623B));
AND2_X1 U_g5500B (.ZN(g5500B),.A2(g4281B),.A1(g1657B));
AND2_X1 U_g2496B (.ZN(g2496B),.A2(g369B),.A1(g374B));
AND2_X1 U_g6756B (.ZN(g6756B),.A2(g5877B),.A1(g3010B));
AND3_X1 U_g8972B (.ZN(g8972B),.A3(FE_OFN73_g8858B),.A2(FE_OFN281_g2216B),.A1(g8085B));
AND2_X1 U_g6622B (.ZN(g6622B),.A2(g6165B),.A1(g336B));
AND2_X1 U_g11639B (.ZN(g11639B),.A2(g7897B),.A1(g11612B));
AND2_X1 U_g9366B (.ZN(g9366B),.A2(FE_OFN53_g9173B),.A1(g1311B));
AND2_X1 U_g11230B (.ZN(g11230B),.A2(g11060B),.A1(g471B));
AND2_X1 U_g10328B (.ZN(g10328B),.A2(FE_OFN269_g109B),.A1(I15507B));
AND2_X1 U_g5024B (.ZN(g5024B),.A2(FE_OFN303_g4678B),.A1(g1284B));
AND2_X1 U_g4364B (.ZN(g4364B),.A2(g4679B),.A1(g1215B));
AND2_X1 U_g9649B (.ZN(g9649B),.A2(g9205B),.A1(g916B));
AND2_X1 U_g5795B (.ZN(g5795B),.A2(g5261B),.A1(g1543B));
AND2_X1 U_g5737B (.ZN(g5737B),.A2(FE_OFN321_g5261B),.A1(g1524B));
AND2_X1 U_g6841B (.ZN(g6841B),.A2(FE_OFN180_g5354B),.A1(g1400B));
AND2_X1 U_g4054B (.ZN(g4054B),.A2(g2774B),.A1(g1753B));
AND2_X1 U_g6345B (.ZN(g6345B),.A2(FE_OFN346_g4381B),.A1(g5823B));
AND2_X1 U_g11391B (.ZN(g11391B),.A2(g7914B),.A1(g11275B));
AND2_X1 U_g9851B (.ZN(g9851B),.A2(g9764B),.A1(g296B));
AND2_X1 U_g6763B (.ZN(g6763B),.A2(g4381B),.A1(g5802B));
AND2_X1 U_g4770B (.ZN(g4770B),.A2(FE_OFN300_g4002B),.A1(g416B));
AND3_X1 U_I16142B (.ZN(I16142B),.A3(g10507B),.A2(g10509B),.A1(g10511B));
AND2_X1 U_g9698B (.ZN(g9698B),.A2(FE_OFN63_g9474B),.A1(g1571B));
AND2_X1 U_g4725B (.ZN(g4725B),.A2(FE_OFN347_g3914B),.A1(g1032B));
AND2_X1 U_g5477B (.ZN(g5477B),.A2(FE_OFN333_g4294B),.A1(g1887B));
AND2_X1 U_g9964B (.ZN(g9964B),.A2(g9536B),.A1(g9954B));
AND2_X1 U_g5523B (.ZN(g5523B),.A2(g4290B),.A1(g1663B));
AND2_X1 U_g4553B (.ZN(g4553B),.A2(g4002B),.A1(g435B));
AND2_X1 U_g8550B (.ZN(g8550B),.A2(FE_OFN330_g7638B),.A1(g8402B));
AND2_X1 U_g8845B (.ZN(g8845B),.A2(FE_OFN328_g8709B),.A1(g8611B));
AND2_X1 U_g2081B (.ZN(g2081B),.A2(g928B),.A1(g932B));
AND2_X1 U_g6359B (.ZN(g6359B),.A2(FE_OFN320_g5361B),.A1(g281B));
AND2_X1 U_g11586B (.ZN(g11586B),.A2(g11539B),.A1(g1324B));
AND2_X1 U_g11007B (.ZN(g11007B),.A2(FE_OFN13_g10702B),.A1(g5147B));
AND2_X1 U_g5104B (.ZN(g5104B),.A2(g4608B),.A1(g1796B));
AND2_X1 U_g5099B (.ZN(g5099B),.A2(FE_OFN141_g3829B),.A1(g4821B));
AND2_X1 U_g6757B (.ZN(g6757B),.A2(g5919B),.A1(g143B));
AND2_X1 U_g5499B (.ZN(g5499B),.A2(g4679B),.A1(g1627B));
AND2_X1 U_g4389B (.ZN(g4389B),.A2(g3092B),.A1(g3529B));
AND2_X1 U_g6416B (.ZN(g6416B),.A2(FE_OFN217_g5013B),.A1(g3497B));
AND2_X1 U_g9720B (.ZN(g9720B),.A2(g9490B),.A1(g1546B));
AND2_X1 U_g4990B (.ZN(g4990B),.A2(FE_OFN147_g4682B),.A1(g1444B));
AND2_X1 U_g9619B (.ZN(g9619B),.A2(g9010B),.A1(g940B));
AND4_X1 U_I6630B (.ZN(I6630B),.A4(FE_OFN253_g1786B),.A3(FE_OFN236_g1776B),.A2(FE_OFN247_g1771B),.A1(g2677B));
AND2_X1 U_g6047B (.ZN(g6047B),.A2(g4977B),.A1(g2017B));
AND2_X1 U_g9652B (.ZN(g9652B),.A2(FE_OFN39_g9223B),.A1(g953B));
AND3_X1 U_g10515B (.ZN(g10515B),.A3(I16142B),.A2(g10469B),.A1(g10505B));
AND2_X1 U_g9843B (.ZN(g9843B),.A2(g9519B),.A1(g9711B));
AND2_X1 U_g5273B (.ZN(g5273B),.A2(g4776B),.A1(g1074B));
AND2_X1 U_g11465B (.ZN(g11465B),.A2(FE_OFN100_g4421B),.A1(g11232B));
AND2_X1 U_g5044B (.ZN(g5044B),.A2(g1918B),.A1(g4348B));
AND2_X1 U_g11237B (.ZN(g11237B),.A2(g11111B),.A1(g4548B));
AND2_X1 U_g9834B (.ZN(g9834B),.A2(FE_OFN34_g9785B),.A1(g9731B));
AND2_X1 U_g6654B (.ZN(g6654B),.A2(FE_OFN282_g6165B),.A1(g363B));
AND2_X1 U_g5444B (.ZN(g5444B),.A2(FE_OFN290_g4880B),.A1(g1041B));
AND2_X1 U_g3714B (.ZN(g3714B),.A2(g2299B),.A1(g1690B));
AND2_X1 U_g11340B (.ZN(g11340B),.A2(g4285B),.A1(g11285B));
AND2_X1 U_g9598B (.ZN(g9598B),.A2(g9274B),.A1(g119B));
AND2_X1 U_g8097B (.ZN(g8097B),.A2(g7852B),.A1(g5477B));
AND2_X1 U_g8726B (.ZN(g8726B),.A2(g7913B),.A1(g8221B));
AND2_X1 U_g6880B (.ZN(g6880B),.A2(g6557B),.A1(g4816B));
AND2_X1 U_g4338B (.ZN(g4338B),.A2(FE_OFN351_g3913B),.A1(g1157B));
AND2_X1 U_g5543B (.ZN(g5543B),.A2(FE_OFN322_g4449B),.A1(g2979B));
AND3_X1 U_g8960B (.ZN(g8960B),.A3(g8828B),.A2(FE_OFN95_g2216B),.A1(g8085B));
AND2_X1 U_g4109B (.ZN(g4109B),.A2(g3287B),.A1(g806B));
AND2_X1 U_g10759B (.ZN(g10759B),.A2(g10556B),.A1(g10557B));
AND2_X1 U_g9938B (.ZN(g9938B),.A2(FE_OFN67_g9367B),.A1(g9917B));
AND2_X1 U_g10758B (.ZN(g10758B),.A2(FE_OFN293_g3015B),.A1(g10652B));
AND2_X1 U_g4759B (.ZN(g4759B),.A2(FE_OFN300_g4002B),.A1(g406B));
AND2_X1 U_g9909B (.ZN(g9909B),.A2(FE_OFN33_g9454B),.A1(g9891B));
AND2_X1 U_g7127B (.ZN(g7127B),.A2(g2241B),.A1(g6663B));
AND2_X1 U_g11165B (.ZN(g11165B),.A2(FE_OFN13_g10702B),.A1(g476B));
AND2_X1 U_g6234B (.ZN(g6234B),.A2(FE_OFN306_g5128B),.A1(g1424B));
AND2_X1 U_g6328B (.ZN(g6328B),.A2(FE_OFN115_g4807B),.A1(g1260B));
AND2_X1 U_g8401B (.ZN(g8401B),.A2(g8146B),.A1(g677B));
AND2_X1 U_g11006B (.ZN(g11006B),.A2(FE_OFN18_g10702B),.A1(g5125B));
AND2_X1 U_g4865B (.ZN(g4865B),.A2(FE_OFN297_g3015B),.A1(g1080B));
AND2_X1 U_g4715B (.ZN(g4715B),.A2(FE_OFN297_g3015B),.A1(g1077B));
AND3_X1 U_g4604B (.ZN(g4604B),.A3(g2325B),.A2(g3753B),.A1(g3056B));
AND2_X1 U_g5513B (.ZN(g5513B),.A2(g3906B),.A1(g1675B));
AND2_X1 U_g11222B (.ZN(g11222B),.A2(FE_OFN279_g11157B),.A1(g965B));
AND2_X1 U_g4498B (.ZN(g4498B),.A2(FE_OFN302_g3913B),.A1(g1145B));
AND2_X1 U_g6554B (.ZN(g6554B),.A2(g5808B),.A1(g96B));
AND2_X1 U_g7732B (.ZN(g7732B),.A2(FE_OFN226_g3880B),.A1(g5803B));
AND2_X1 U_g9586B (.ZN(g9586B),.A2(FE_OFN53_g9173B),.A1(g1346B));
AND3_X1 U_g5178B (.ZN(g5178B),.A3(g4104B),.A2(FE_OFN223_g4401B),.A1(g2047B));
AND2_X1 U_g4584B (.ZN(g4584B),.A2(g1857B),.A1(g3710B));
AND2_X1 U_g7472B (.ZN(g7472B),.A2(g61B),.A1(FE_OFN83_g2176B));
AND2_X1 U_g11253B (.ZN(g11253B),.A2(g11083B),.A1(g981B));
AND2_X1 U_g5182B (.ZN(g5182B),.A2(FE_OFN303_g4678B),.A1(g1240B));
AND2_X1 U_g9860B (.ZN(g9860B),.A2(g9778B),.A1(g1598B));
AND2_X1 U_g11600B (.ZN(g11600B),.A2(g11575B),.A1(g1346B));
AND2_X1 U_g9710B (.ZN(g9710B),.A2(FE_OFN63_g9474B),.A1(g1586B));
AND2_X1 U_g9645B (.ZN(g9645B),.A2(FE_OFN51_g9111B),.A1(g1203B));
AND2_X1 U_g11236B (.ZN(g11236B),.A2(g11111B),.A1(g4537B));
AND2_X1 U_g4162B (.ZN(g4162B),.A2(g1845B),.A1(g3106B));
AND2_X1 U_g6090B (.ZN(g6090B),.A2(g5627B),.A1(g553B));
AND2_X1 U_g9691B (.ZN(g9691B),.A2(g9432B),.A1(g269B));
AND2_X1 U_g11372B (.ZN(g11372B),.A2(g4285B),.A1(g11316B));
AND2_X1 U_g6823B (.ZN(g6823B),.A2(g5354B),.A1(g1368B));
AND2_X1 U_g11175B (.ZN(g11175B),.A2(FE_OFN20_g10702B),.A1(g501B));
AND2_X1 U_g8068B (.ZN(g8068B),.A2(FE_OFN198_g7697B),.A1(g664B));
AND2_X1 U_g9607B (.ZN(g9607B),.A2(g9274B),.A1(g12B));
AND2_X1 U_g9962B (.ZN(g9962B),.A2(FE_OFN280_g9536B),.A1(g9952B));
AND2_X1 U_g6348B (.ZN(g6348B),.A2(FE_OFN320_g5361B),.A1(g296B));
AND2_X1 U_g9659B (.ZN(g9659B),.A2(FE_OFN39_g9223B),.A1(g956B));
AND2_X1 U_g9358B (.ZN(g9358B),.A2(FE_OFN47_g9151B),.A1(g1318B));
AND2_X1 U_g3104B (.ZN(g3104B),.A2(I6317B),.A1(I6316B));
AND2_X1 U_g4486B (.ZN(g4486B),.A2(g4679B),.A1(g1711B));
AND2_X1 U_g9587B (.ZN(g9587B),.A2(g8995B),.A1(g892B));
AND2_X1 U_g5632B (.ZN(g5632B),.A2(I5435B),.A1(g1636B));
AND2_X4 U_g9111B (.ZN(g9111B),.A2(FE_OFN276_g48B),.A1(g8965B));
AND2_X1 U_g4881B (.ZN(g4881B),.A2(FE_OFN347_g3914B),.A1(g991B));
AND2_X1 U_g11209B (.ZN(g11209B),.A2(FE_OFN79_g8700B),.A1(g10712B));
AND2_X1 U_g8848B (.ZN(g8848B),.A2(FE_OFN328_g8709B),.A1(g8715B));
AND2_X1 U_g4070B (.ZN(g4070B),.A2(g2330B),.A1(g3263B));
AND2_X1 U_g6463B (.ZN(g6463B),.A2(I9237B),.A1(FE_OFN277_g48B));
AND4_X1 U_I5689B (.ZN(I5689B),.A4(g1432B),.A3(g1428B),.A2(g1424B),.A1(g1419B));
AND2_X1 U_g7820B (.ZN(g7820B),.A2(FE_OFN209_g6863B),.A1(g1896B));
AND2_X1 U_g11021B (.ZN(g11021B),.A2(FE_OFN7_g10702B),.A1(g448B));
AND2_X1 U_g5917B (.ZN(g5917B),.A2(g85B),.A1(g1044B));
AND2_X1 U_g6619B (.ZN(g6619B),.A2(FE_OFN97_I8869B),.A1(g49B));
AND2_X1 U_g6318B (.ZN(g6318B),.A2(FE_OFN118_g4807B),.A1(g1300B));
AND2_X1 U_g6872B (.ZN(g6872B),.A2(FE_OFN213_g6003B),.A1(g1896B));
AND2_X1 U_g11320B (.ZN(g11320B),.A2(g4379B),.A1(g11201B));
AND2_X1 U_g10514B (.ZN(g10514B),.A2(FE_OFN370_g4525B),.A1(g10489B));
AND2_X1 U_g4006B (.ZN(g4006B),.A2(FE_OFN266_g18B),.A1(g201B));
AND2_X1 U_g9853B (.ZN(g9853B),.A2(g9764B),.A1(g299B));
AND2_X1 U_g11274B (.ZN(g11274B),.A2(g11199B),.A1(g4771B));
AND2_X1 U_g6193B (.ZN(g6193B),.A2(FE_OFN306_g5128B),.A1(g1419B));
AND2_X1 U_g8119B (.ZN(g8119B),.A2(FE_OFN207_g6863B),.A1(g5526B));
AND2_X1 U_g9420B (.ZN(g9420B),.A2(FE_OFN50_g9030B),.A1(g1747B));
AND2_X1 U_g5233B (.ZN(g5233B),.A2(g4492B),.A1(FE_OFN252_g1791B));
AND2_X1 U_g7581B (.ZN(g7581B),.A2(g5420B),.A1(g7092B));
AND2_X1 U_g6549B (.ZN(g6549B),.A2(g5808B),.A1(g95B));
AND2_X1 U_g11464B (.ZN(g11464B),.A2(FE_OFN100_g4421B),.A1(g11231B));
AND2_X1 U_g4801B (.ZN(g4801B),.A2(FE_OFN307_g4010B),.A1(g516B));
AND2_X1 U_g6834B (.ZN(g6834B),.A2(FE_OFN178_g5354B),.A1(g1365B));
AND2_X1 U_g4487B (.ZN(g4487B),.A2(g3906B),.A1(g1718B));
AND2_X1 U_g2939B (.ZN(g2939B),.A2(g1687B),.A1(FE_OFN241_g1690B));
AND2_X1 U_g7060B (.ZN(g7060B),.A2(g5521B),.A1(g6739B));
AND2_X1 U_g5770B (.ZN(g5770B),.A2(g5128B),.A1(g3585B));
AND2_X1 U_g5725B (.ZN(g5725B),.A2(FE_OFN353_g5117B),.A1(g1580B));
AND2_X1 U_g11641B (.ZN(g11641B),.A2(g7897B),.A1(g11615B));
AND2_X1 U_g2544B (.ZN(g2544B),.A2(g1336B),.A1(g1341B));
AND2_X1 U_g11292B (.ZN(g11292B),.A2(g4379B),.A1(g11252B));
AND2_X1 U_g5532B (.ZN(g5532B),.A2(g4273B),.A1(g1681B));
AND2_X1 U_g11153B (.ZN(g11153B),.A2(g10788B),.A1(g3771B));
AND2_X1 U_g9905B (.ZN(g9905B),.A2(g9680B),.A1(g9872B));
AND2_X1 U_g7739B (.ZN(g7739B),.A2(g3880B),.A1(g5820B));
AND2_X1 U_g6321B (.ZN(g6321B),.A2(FE_OFN118_g4807B),.A1(g1284B));
AND2_X1 U_g8386B (.ZN(g8386B),.A2(g8220B),.A1(g5257B));
AND3_X1 U_g8975B (.ZN(g8975B),.A3(FE_OFN73_g8858B),.A2(FE_OFN281_g2216B),.A1(g8089B));
AND2_X1 U_g2306B (.ZN(g2306B),.A2(g1218B),.A1(g1223B));
AND2_X1 U_g6625B (.ZN(g6625B),.A2(g6081B),.A1(g1218B));
AND2_X1 U_g7937B (.ZN(g7937B),.A2(FE_OFN292_g3015B),.A1(g5274B));
AND2_X2 U_g10788B (.ZN(g10788B),.A2(g10702B),.A1(g8303B));
AND2_X1 U_g10325B (.ZN(g10325B),.A2(FE_OFN352_g109B),.A1(I15503B));
AND2_X1 U_g8170B (.ZN(g8170B),.A2(FE_OFN89_I11360B),.A1(g36B));
AND2_X1 U_g5706B (.ZN(g5706B),.A2(FE_OFN315_g5117B),.A1(g1574B));
AND2_X1 U_g2756B (.ZN(g2756B),.A2(g2081B),.A1(g936B));
AND2_X1 U_g8821B (.ZN(g8821B),.A2(FE_OFN328_g8709B),.A1(g8643B));
AND2_X1 U_g10946B (.ZN(g10946B),.A2(FE_OFN9_g10702B),.A1(g5225B));
AND2_X1 U_g4169B (.ZN(g4169B),.A2(g3060B),.A1(FE_OFN237_g1806B));
AND2_X1 U_g5029B (.ZN(g5029B),.A2(FE_OFN288_g4263B),.A1(g1077B));
AND2_X1 U_g11164B (.ZN(g11164B),.A2(FE_OFN13_g10702B),.A1(g3513B));
AND2_X1 U_g4007B (.ZN(g4007B),.A2(g2276B),.A1(FE_OFN247_g1771B));
AND2_X1 U_g4059B (.ZN(g4059B),.A2(g2774B),.A1(g1756B));
AND2_X1 U_g4868B (.ZN(g4868B),.A2(FE_OFN347_g3914B),.A1(g1027B));
AND2_X1 U_g5675B (.ZN(g5675B),.A2(FE_OFN365_g5361B),.A1(g131B));
AND2_X1 U_g4718B (.ZN(g4718B),.A2(g3943B),.A1(g650B));
AND2_X1 U_g10682B (.ZN(g10682B),.A2(FE_OFN136_g3863B),.A1(g10381B));
AND2_X1 U_g6687B (.ZN(g6687B),.A2(I9326B),.A1(g92B));
AND2_X1 U_g7704B (.ZN(g7704B),.A2(FE_OFN191_g6488B),.A1(g682B));
AND2_X1 U_g4582B (.ZN(g4582B),.A2(g4010B),.A1(g525B));
AND2_X1 U_g4261B (.ZN(g4261B),.A2(FE_OFN347_g3914B),.A1(g1019B));
AND2_X1 U_g3422B (.ZN(g3422B),.A2(FE_OFN324_g18B),.A1(g225B));
AND2_X1 U_g5745B (.ZN(g5745B),.A2(FE_OFN321_g5261B),.A1(g1549B));
AND2_X1 U_g8387B (.ZN(g8387B),.A2(g8220B),.A1(g5258B));
AND2_X1 U_g7954B (.ZN(g7954B),.A2(g7512B),.A1(g49B));
AND2_X1 U_g11283B (.ZN(g11283B),.A2(g11239B),.A1(g4804B));
AND2_X1 U_g8461B (.ZN(g8461B),.A2(FE_OFN210_g7246B),.A1(g8298B));
AND2_X1 U_g10760B (.ZN(g10760B),.A2(g10554B),.A1(g10555B));
AND2_X1 U_g11492B (.ZN(g11492B),.A2(g4807B),.A1(g11480B));
AND3_X1 U_g7032B (.ZN(g7032B),.A3(I7048B),.A2(g6626B),.A1(g109B));
AND2_X4 U_g9151B (.ZN(g9151B),.A2(FE_OFN276_g48B),.A1(g8967B));
AND2_X1 U_g6341B (.ZN(g6341B),.A2(FE_OFN319_g5361B),.A1(g272B));
AND2_X1 U_g10506B (.ZN(g10506B),.A2(FE_OFN241_g1690B),.A1(g10007B));
AND2_X1 U_g9648B (.ZN(g9648B),.A2(FE_OFN62_g9274B),.A1(g16B));
AND2_X1 U_g7453B (.ZN(g7453B),.A2(g52B),.A1(FE_OFN86_g2176B));
AND2_X1 U_g6525B (.ZN(g6525B),.A2(FE_OFN343_I5565B),.A1(g5995B));
AND2_X1 U_g6645B (.ZN(g6645B),.A2(FE_OFN97_I8869B),.A1(g67B));
AND2_X1 U_g5707B (.ZN(g5707B),.A2(FE_OFN353_g5117B),.A1(g1595B));
AND2_X1 U_g8046B (.ZN(g8046B),.A2(FE_OFN305_g5151B),.A1(g7548B));
AND2_X1 U_g11091B (.ZN(g11091B),.A2(FE_OFN4_g10950B),.A1(g833B));
AND2_X1 U_g11174B (.ZN(g11174B),.A2(FE_OFN21_g10702B),.A1(g496B));
AND2_X4 U_g9010B (.ZN(g9010B),.A2(g8930B),.A1(FE_OFN277_g48B));
AND2_X1 U_g8403B (.ZN(g8403B),.A2(g8220B),.A1(g5276B));
AND2_X1 U_g5201B (.ZN(g5201B),.A2(g4678B),.A1(g1250B));
AND2_X1 U_g8841B (.ZN(g8841B),.A2(FE_OFN328_g8709B),.A1(g8605B));
AND2_X1 U_g6879B (.ZN(g6879B),.A2(FE_OFN213_g6003B),.A1(g1914B));
AND2_X2 U_g8763B (.ZN(g8763B),.A2(g8451B),.A1(I9880B));
AND2_X1 U_g4502B (.ZN(g4502B),.A2(g3938B),.A1(g2031B));
AND2_X1 U_g9839B (.ZN(g9839B),.A2(g9747B),.A1(g9702B));
AND2_X1 U_g6358B (.ZN(g6358B),.A2(FE_OFN346_g4381B),.A1(g5841B));
AND2_X1 U_g5575B (.ZN(g5575B),.A2(FE_OFN367_g3521B),.A1(g1618B));
AND2_X1 U_g4940B (.ZN(g4940B),.A2(FE_OFN310_g4336B),.A1(g1984B));
AND2_X1 U_g8107B (.ZN(g8107B),.A2(g7852B),.A1(g5502B));
AND2_X1 U_g10240B (.ZN(g10240B),.A2(g9082B),.A1(g9974B));
AND2_X1 U_g11192B (.ZN(g11192B),.A2(g10927B),.A1(g4759B));
AND2_X1 U_g9618B (.ZN(g9618B),.A2(g9205B),.A1(g910B));
AND2_X1 U_g5539B (.ZN(g5539B),.A2(g4273B),.A1(g1684B));
AND2_X1 U_g8416B (.ZN(g8416B),.A2(FE_OFN187_g7638B),.A1(g731B));
AND2_X1 U_g9693B (.ZN(g9693B),.A2(FE_OFN59_g9432B),.A1(g275B));
AND2_X1 U_g11553B (.ZN(g11553B),.A2(g11519B),.A1(g1771B));
AND2_X1 U_g8047B (.ZN(g8047B),.A2(FE_OFN177_g5919B),.A1(g7557B));
AND2_X1 U_g5268B (.ZN(g5268B),.A2(g4263B),.A1(g1098B));
AND2_X1 U_g9555B (.ZN(g9555B),.A2(FE_OFN325_g18B),.A1(g9107B));
AND2_X1 U_g6180B (.ZN(g6180B),.A2(g5128B),.A1(g1453B));
AND2_X1 U_g6832B (.ZN(g6832B),.A2(FE_OFN179_g5354B),.A1(g1383B));
AND2_X1 U_g10633B (.ZN(g10633B),.A2(g3829B),.A1(g10381B));
AND2_X1 U_g7894B (.ZN(g7894B),.A2(FE_OFN366_g3521B),.A1(g5317B));
AND2_X1 U_g8654B (.ZN(g8654B),.A2(FE_OFN348_g3015B),.A1(g8266B));
AND2_X1 U_g9621B (.ZN(g9621B),.A2(FE_OFN46_g9125B),.A1(g1179B));
AND2_X1 U_g6794B (.ZN(g6794B),.A2(FE_OFN346_g4381B),.A1(g5819B));
AND2_X1 U_g9313B (.ZN(g9313B),.A2(FE_OFN275_g48B),.A1(g8876B));
AND2_X1 U_g3412B (.ZN(g3412B),.A2(g18B),.A1(g219B));
AND2_X1 U_g7661B (.ZN(g7661B),.A2(g2251B),.A1(g7127B));
AND3_X1 U_g2800B (.ZN(g2800B),.A3(g591B),.A2(g2369B),.A1(g2399B));
AND2_X1 U_g3706B (.ZN(g3706B),.A2(g3268B),.A1(g471B));
AND2_X1 U_g9908B (.ZN(g9908B),.A2(FE_OFN33_g9454B),.A1(g9760B));
AND2_X1 U_g3429B (.ZN(g3429B),.A2(g18B),.A1(g231B));
AND2_X1 U_g6628B (.ZN(g6628B),.A2(FE_OFN282_g6165B),.A1(g351B));
AND2_X1 U_g5470B (.ZN(g5470B),.A2(g4880B),.A1(g1044B));
AND2_X1 U_g7526B (.ZN(g7526B),.A2(g73B),.A1(FE_OFN87_g2176B));
AND2_X1 U_g5897B (.ZN(g5897B),.A2(g5354B),.A1(g2204B));
AND2_X1 U_g5025B (.ZN(g5025B),.A2(FE_OFN153_g4640B),.A1(g1482B));
AND2_X1 U_g6204B (.ZN(g6204B),.A2(FE_OFN200_g4921B),.A1(g3738B));
AND2_X1 U_g4048B (.ZN(g4048B),.A2(g2774B),.A1(g1750B));
AND3_X1 U_g8935B (.ZN(g8935B),.A3(g8849B),.A2(FE_OFN95_g2216B),.A1(g8106B));
AND2_X1 U_g3281B (.ZN(g3281B),.A2(g2525B),.A1(g766B));
AND2_X1 U_g9593B (.ZN(g9593B),.A2(FE_OFN42_g9205B),.A1(g898B));
AND2_X1 U_g4827B (.ZN(g4827B),.A2(FE_OFN324_g18B),.A1(g213B));
AND2_X1 U_g10701B (.ZN(g10701B),.A2(g10500B),.A1(g10501B));
AND2_X1 U_g10777B (.ZN(g10777B),.A2(g3015B),.A1(g10733B));
AND2_X1 U_g8130B (.ZN(g8130B),.A2(g7952B),.A1(g1936B));
AND2_X1 U_g9965B (.ZN(g9965B),.A2(FE_OFN280_g9536B),.A1(g9955B));
AND2_X1 U_g3684B (.ZN(g3684B),.A2(g3015B),.A1(g1710B));
AND2_X1 U_g11213B (.ZN(g11213B),.A2(FE_OFN279_g11157B),.A1(g947B));
AND2_X1 U_g5006B (.ZN(g5006B),.A2(FE_OFN154_g4640B),.A1(g1462B));
AND2_X1 U_g9933B (.ZN(g9933B),.A2(g9624B),.A1(g9912B));
AND2_X1 U_g8554B (.ZN(g8554B),.A2(FE_OFN330_g7638B),.A1(g8407B));
AND2_X1 U_g9641B (.ZN(g9641B),.A2(g9205B),.A1(g913B));
AND2_X1 U_g6123B (.ZN(g6123B),.A2(FE_OFN310_g4336B),.A1(g3662B));
AND2_X1 U_g6323B (.ZN(g6323B),.A2(FE_OFN116_g4807B),.A1(g1235B));
AND2_X1 U_g10766B (.ZN(g10766B),.A2(FE_OFN131_g3015B),.A1(g10646B));
AND2_X1 U_g6666B (.ZN(g6666B),.A2(g5836B),.A1(g89B));
AND2_X1 U_g4994B (.ZN(g4994B),.A2(FE_OFN154_g4640B),.A1(g1504B));
AND2_X1 U_g5755B (.ZN(g5755B),.A2(FE_OFN179_g5354B),.A1(g5103B));
AND2_X1 U_g11592B (.ZN(g11592B),.A2(g11561B),.A1(g3717B));
AND2_X1 U_g6351B (.ZN(g6351B),.A2(g48B),.A1(I9237B));
AND2_X1 U_g6875B (.ZN(g6875B),.A2(FE_OFN213_g6003B),.A1(g1905B));
AND2_X1 U_g4816B (.ZN(g4816B),.A2(g2336B),.A1(g4070B));
AND2_X1 U_g9658B (.ZN(g9658B),.A2(g9240B),.A1(g947B));
AND2_X1 U_g6530B (.ZN(g6530B),.A2(FE_OFN141_g3829B),.A1(g6207B));
AND2_X1 U_g8366B (.ZN(g8366B),.A2(g7265B),.A1(g8199B));
AND2_X1 U_g9835B (.ZN(g9835B),.A2(FE_OFN34_g9785B),.A1(g9735B));
AND2_X1 U_g6655B (.ZN(g6655B),.A2(I9326B),.A1(g88B));
AND3_X1 U_g5445B (.ZN(g5445B),.A3(g109B),.A2(g3875B),.A1(FE_OFN184_I7048B));
AND2_X1 U_g5173B (.ZN(g5173B),.A2(g4671B),.A1(g1110B));
AND2_X1 U_g7970B (.ZN(g7970B),.A2(g7438B),.A1(g7384B));
AND2_X1 U_g3098B (.ZN(g3098B),.A2(g2198B),.A1(g2331B));
AND2_X1 U_g5491B (.ZN(g5491B),.A2(g4289B),.A1(g1624B));
AND2_X1 U_g9271B (.ZN(g9271B),.A2(g8949B),.A1(g6109B));
AND2_X1 U_g11152B (.ZN(g11152B),.A2(g10883B),.A1(g369B));
AND2_X1 U_g9611B (.ZN(g9611B),.A2(g9010B),.A1(g936B));
AND2_X1 U_g6410B (.ZN(g6410B),.A2(FE_OFN217_g5013B),.A1(g2804B));
AND2_X1 U_g10451B (.ZN(g10451B),.A2(g2024B),.A1(g10444B));
AND2_X1 U_g4397B (.ZN(g4397B),.A2(g639B),.A1(g3475B));
AND2_X1 U_g7224B (.ZN(g7224B),.A2(g6447B),.A1(g5398B));
AND2_X1 U_g5602B (.ZN(g5602B),.A2(FE_OFN357_g3521B),.A1(g1624B));
AND2_X2 U_g4421B (.ZN(g4421B),.A2(g750B),.A1(g2057B));
AND2_X1 U_g6884B (.ZN(g6884B),.A2(g6557B),.A1(g5569B));
AND2_X1 U_g6839B (.ZN(g6839B),.A2(FE_OFN180_g5354B),.A1(g1397B));
AND3_X1 U_g8964B (.ZN(g8964B),.A3(g8849B),.A2(FE_OFN92_g2216B),.A1(g8255B));
AND2_X1 U_g8260B (.ZN(g8260B),.A2(g7907B),.A1(g940B));
AND2_X1 U_g11413B (.ZN(g11413B),.A2(g10679B),.A1(g11217B));
AND2_X1 U_g4950B (.ZN(g4950B),.A2(FE_OFN146_g4682B),.A1(g1415B));
AND2_X1 U_g5535B (.ZN(g5535B),.A2(FE_OFN366_g3521B),.A1(g572B));
AND2_X1 U_g7277B (.ZN(g7277B),.A2(g731B),.A1(g6772B));
AND2_X1 U_g8463B (.ZN(g8463B),.A2(FE_OFN211_g7246B),.A1(g8301B));
AND2_X1 U_g3268B (.ZN(g3268B),.A2(g2511B),.A1(FE_OFN248_g466B));
AND2_X1 U_g10785B (.ZN(g10785B),.A2(g4467B),.A1(g10728B));
AND2_X1 U_g6618B (.ZN(g6618B),.A2(FE_OFN219_g5557B),.A1(g658B));
AND2_X1 U_g6235B (.ZN(g6235B),.A2(g5613B),.A1(g569B));
AND2_X1 U_g10950B (.ZN(g10950B),.A2(g6355B),.A1(g10788B));
AND2_X1 U_g4723B (.ZN(g4723B),.A2(g627B),.A1(g3626B));
AND2_X1 U_g8720B (.ZN(g8720B),.A2(g7905B),.A1(g8206B));
AND2_X1 U_g6693B (.ZN(g6693B),.A2(I9326B),.A1(g93B));
AND2_X1 U_g11020B (.ZN(g11020B),.A2(FE_OFN7_g10702B),.A1(g452B));
AND2_X1 U_g11583B (.ZN(g11583B),.A2(g11539B),.A1(g1314B));
AND2_X1 U_g8118B (.ZN(g8118B),.A2(g7949B),.A1(g1900B));
AND2_X1 U_g8167B (.ZN(g8167B),.A2(FE_OFN89_I11360B),.A1(g33B));
AND2_X1 U_g6334B (.ZN(g6334B),.A2(FE_OFN180_g5354B),.A1(g1389B));
AND2_X1 U_g7892B (.ZN(g7892B),.A2(g3814B),.A1(g5308B));
AND2_X1 U_g8652B (.ZN(g8652B),.A2(FE_OFN119_g3015B),.A1(g8264B));
AND2_X1 U_g5721B (.ZN(g5721B),.A2(FE_OFN353_g5117B),.A1(g1577B));
AND2_X1 U_g10367B (.ZN(g10367B),.A2(FE_OFN234_g2024B),.A1(g10362B));
AND2_X1 U_g9901B (.ZN(g9901B),.A2(FE_OFN69_g9392B),.A1(g9719B));
AND2_X1 U_g6792B (.ZN(g6792B),.A2(FE_OFN319_g5361B),.A1(g290B));
AND2_X1 U_g11282B (.ZN(g11282B),.A2(g11203B),.A1(g4801B));
AND2_X1 U_g7945B (.ZN(g7945B),.A2(g7473B),.A1(g67B));
AND3_X1 U_g8971B (.ZN(g8971B),.A3(FE_OFN73_g8858B),.A2(FE_OFN281_g2216B),.A1(g8081B));
AND2_X1 U_g11302B (.ZN(g11302B),.A2(g11243B),.A1(g4582B));
AND2_X1 U_g4585B (.ZN(g4585B),.A2(g4010B),.A1(g521B));
AND2_X1 U_g6621B (.ZN(g6621B),.A2(I8869B),.A1(g52B));
AND2_X1 U_g5502B (.ZN(g5502B),.A2(FE_OFN333_g4294B),.A1(g1932B));
AND2_X1 U_g11105B (.ZN(g11105B),.A2(g10937B),.A1(g3634B));
AND2_X1 U_g7709B (.ZN(g7709B),.A2(FE_OFN322_g4449B),.A1(g5942B));
AND2_X1 U_g8598B (.ZN(g8598B),.A2(FE_OFN210_g7246B),.A1(g8471B));
AND2_X1 U_g7140B (.ZN(g7140B),.A2(g6716B),.A1(g5221B));
AND2_X1 U_g9600B (.ZN(g9600B),.A2(FE_OFN42_g9205B),.A1(g904B));
AND2_X1 U_g9864B (.ZN(g9864B),.A2(g9778B),.A1(g1604B));
AND2_X1 U_g11640B (.ZN(g11640B),.A2(g7897B),.A1(g11613B));
AND2_X1 U_g5188B (.ZN(g5188B),.A2(g794B),.A1(g798B));
AND2_X1 U_g7435B (.ZN(g7435B),.A2(g6403B),.A1(g7260B));
AND2_X1 U_g7876B (.ZN(g7876B),.A2(FE_OFN366_g3521B),.A1(g5278B));
AND2_X1 U_g5030B (.ZN(g5030B),.A2(FE_OFN303_g4678B),.A1(g1280B));
AND2_X1 U_g4058B (.ZN(g4058B),.A2(FE_OFN224_g2276B),.A1(FE_OFN252_g1791B));
AND2_X1 U_g6776B (.ZN(g6776B),.A2(FE_OFN111_g3914B),.A1(g5809B));
AND2_X1 U_g4890B (.ZN(g4890B),.A2(g4739B),.A1(g630B));
AND2_X1 U_g2525B (.ZN(g2525B),.A2(g758B),.A1(g762B));
AND2_X1 U_g10301B (.ZN(g10301B),.A2(g10025B),.A1(g8700B));
AND2_X1 U_g4505B (.ZN(g4505B),.A2(FE_OFN287_g3586B),.A1(g354B));
AND2_X1 U_g9623B (.ZN(g9623B),.A2(FE_OFN62_g9274B),.A1(g17B));
AND2_X1 U_g10739B (.ZN(g10739B),.A2(g3368B),.A1(g10676B));
AND2_X1 U_g11027B (.ZN(g11027B),.A2(FE_OFN17_g10702B),.A1(g391B));
AND2_X1 U_g10738B (.ZN(g10738B),.A2(FE_OFN131_g3015B),.A1(g10599B));
AND2_X1 U_g8687B (.ZN(g8687B),.A2(FE_OFN189_g7638B),.A1(g8558B));
AND2_X1 U_g6360B (.ZN(g6360B),.A2(FE_OFN319_g5361B),.A1(g302B));
AND2_X1 U_g9871B (.ZN(g9871B),.A2(g9802B),.A1(g1564B));
AND2_X1 U_g5108B (.ZN(g5108B),.A2(g4608B),.A1(g1801B));
AND2_X1 U_g11248B (.ZN(g11248B),.A2(g11083B),.A1(g976B));
AND2_X1 U_g4992B (.ZN(g4992B),.A2(FE_OFN147_g4682B),.A1(g1407B));
AND2_X1 U_g11552B (.ZN(g11552B),.A2(FE_OFN27_g11519B),.A1(g2677B));
AND2_X1 U_g9651B (.ZN(g9651B),.A2(g9240B),.A1(g944B));
AND2_X1 U_g11204B (.ZN(g11204B),.A2(g11083B),.A1(g971B));
AND2_X1 U_g7824B (.ZN(g7824B),.A2(FE_OFN206_g6863B),.A1(g1932B));
AND2_X1 U_g4480B (.ZN(g4480B),.A2(FE_OFN302_g3913B),.A1(g1133B));
AND2_X1 U_g6179B (.ZN(g6179B),.A2(g5354B),.A1(g5115B));
AND2_X1 U_g7590B (.ZN(g7590B),.A2(g5420B),.A1(g7102B));
AND2_X1 U_g9384B (.ZN(g9384B),.A2(g9223B),.A1(g968B));
AND2_X1 U_g3407B (.ZN(g3407B),.A2(FE_OFN352_g109B),.A1(g2561B));
AND2_X1 U_g9838B (.ZN(g9838B),.A2(g9754B),.A1(g9700B));
AND2_X1 U_g10661B (.ZN(g10661B),.A2(FE_OFN119_g3015B),.A1(g10594B));
AND2_X1 U_g11380B (.ZN(g11380B),.A2(g4285B),.A1(g11321B));
AND3_X1 U_g8879B (.ZN(g8879B),.A3(FE_OFN73_g8858B),.A2(FE_OFN281_g2216B),.A1(g8110B));
AND2_X1 U_g7930B (.ZN(g7930B),.A2(FE_OFN343_I5565B),.A1(g7621B));
AND3_X1 U_g8962B (.ZN(g8962B),.A3(g8828B),.A2(FE_OFN95_g2216B),.A1(g8089B));
AND2_X1 U_g10715B (.ZN(g10715B),.A2(g10584B),.A1(g2272B));
AND2_X1 U_g8659B (.ZN(g8659B),.A2(FE_OFN298_g3015B),.A1(g8269B));
AND2_X4 U_g3015B (.ZN(g3015B),.A2(I6260B),.A1(g2028B));
AND2_X1 U_g9643B (.ZN(g9643B),.A2(FE_OFN39_g9223B),.A1(g950B));
AND2_X4 U_g9205B (.ZN(g9205B),.A2(g8957B),.A1(FE_OFN276_g48B));
AND2_X1 U_g5538B (.ZN(g5538B),.A2(FE_OFN288_g4263B),.A1(g1669B));
AND2_X1 U_g4000B (.ZN(g4000B),.A2(g2774B),.A1(g1744B));
AND2_X1 U_g4126B (.ZN(g4126B),.A2(g3060B),.A1(FE_OFN253_g1786B));
AND2_X1 U_g4400B (.ZN(g4400B),.A2(FE_OFN137_g3829B),.A1(g4088B));
AND2_X1 U_g2794B (.ZN(g2794B),.A2(I5887B),.A1(I5886B));
AND2_X1 U_g4760B (.ZN(g4760B),.A2(FE_OFN307_g4010B),.A1(g486B));
AND2_X1 U_g6238B (.ZN(g6238B),.A2(FE_OFN289_g4679B),.A1(g572B));
AND2_X1 U_g10784B (.ZN(g10784B),.A2(g4467B),.A1(g10727B));
AND2_X1 U_g8174B (.ZN(g8174B),.A2(FE_OFN89_I11360B),.A1(g38B));
AND2_X1 U_g6332B (.ZN(g6332B),.A2(FE_OFN180_g5354B),.A1(g1374B));
AND2_X1 U_g5067B (.ZN(g5067B),.A2(g4811B),.A1(g305B));
AND2_X1 U_g5418B (.ZN(g5418B),.A2(FE_OFN357_g3521B),.A1(g1512B));
AND2_X1 U_g10297B (.ZN(g10297B),.A2(g10001B),.A1(FE_OFN79_g8700B));
AND2_X1 U_g6353B (.ZN(g6353B),.A2(FE_OFN320_g5361B),.A1(g299B));
AND2_X1 U_g11026B (.ZN(g11026B),.A2(FE_OFN14_g10702B),.A1(g386B));
AND2_X1 U_g11212B (.ZN(g11212B),.A2(FE_OFN279_g11157B),.A1(g944B));
AND2_X1 U_g6744B (.ZN(g6744B),.A2(FE_OFN218_g5557B),.A1(g4828B));
AND2_X1 U_g5493B (.ZN(g5493B),.A2(FE_OFN333_g4294B),.A1(g1923B));
AND2_X1 U_g10671B (.ZN(g10671B),.A2(g9473B),.A1(g10411B));
AND2_X1 U_g4383B (.ZN(g4383B),.A2(FE_OFN141_g3829B),.A1(g2517B));
AND2_X1 U_g5256B (.ZN(g5256B),.A2(g627B),.A1(g4297B));
AND2_X1 U_g4220B (.ZN(g4220B),.A2(g3539B),.A1(g105B));
AND2_X1 U_g8380B (.ZN(g8380B),.A2(FE_OFN333_g4294B),.A1(g8252B));
AND2_X1 U_g7071B (.ZN(g7071B),.A2(g6586B),.A1(g5030B));
AND2_X1 U_g4779B (.ZN(g4779B),.A2(FE_OFN307_g4010B),.A1(g501B));
AND2_X1 U_g9613B (.ZN(g9613B),.A2(FE_OFN46_g9125B),.A1(g1176B));
AND2_X1 U_g7705B (.ZN(g7705B),.A2(g4336B),.A1(g5935B));
AND2_X1 U_g9269B (.ZN(g9269B),.A2(FE_OFN266_g18B),.A1(g8933B));
AND2_X1 U_g5181B (.ZN(g5181B),.A2(g802B),.A1(g806B));
AND2_X1 U_g4977B (.ZN(g4977B),.A2(g4807B),.A1(g4567B));
AND2_X1 U_g7948B (.ZN(g7948B),.A2(g7497B),.A1(g70B));
AND2_X1 U_g11149B (.ZN(g11149B),.A2(FE_OFN278_g10927B),.A1(g324B));
AND2_X1 U_g9862B (.ZN(g9862B),.A2(g9778B),.A1(g1601B));
AND2_X1 U_g11387B (.ZN(g11387B),.A2(g3629B),.A1(g11077B));
AND2_X1 U_g7955B (.ZN(g7955B),.A2(g7516B),.A1(g76B));
AND2_X1 U_g4161B (.ZN(g4161B),.A2(g3060B),.A1(FE_OFN251_g1801B));
AND2_X1 U_g11148B (.ZN(g11148B),.A2(g10788B),.A1(g2321B));
AND2_X1 U_g9712B (.ZN(g9712B),.A2(FE_OFN70_g9490B),.A1(g1528B));
AND2_X1 U_g8931B (.ZN(g8931B),.A2(g8164B),.A1(g8642B));
AND2_X1 U_g11097B (.ZN(g11097B),.A2(g10883B),.A1(g378B));
AND3_X1 U_g5421B (.ZN(g5421B),.A3(g3819B),.A2(g109B),.A1(FE_OFN184_I7048B));
AND2_X1 U_g11104B (.ZN(g11104B),.A2(g10937B),.A1(g2963B));
AND2_X1 U_g5263B (.ZN(g5263B),.A2(FE_OFN335_g4737B),.A1(g709B));
AND2_X1 U_g6092B (.ZN(g6092B),.A2(FE_OFN273_g85B),.A1(g1059B));
AND2_X1 U_g4999B (.ZN(g4999B),.A2(FE_OFN154_g4640B),.A1(g1499B));
AND4_X1 U_I6338B (.ZN(I6338B),.A4(g2446B),.A3(g2451B),.A2(g2456B),.A1(g2475B));
AND3_X1 U_g7409B (.ZN(g7409B),.A3(g6858B),.A2(g632B),.A1(g4976B));
AND2_X1 U_g4103B (.ZN(g4103B),.A2(g3060B),.A1(FE_OFN247_g1771B));
AND4_X1 U_I6309B (.ZN(I6309B),.A4(g2475B),.A3(g2456B),.A2(g2451B),.A1(g2446B));
AND2_X1 U_g6580B (.ZN(g6580B),.A2(g5944B),.A1(FE_OFN251_g1801B));
AND2_X1 U_g5631B (.ZN(g5631B),.A2(FE_OFN291_g4880B),.A1(g1056B));
AND2_X1 U_g9414B (.ZN(g9414B),.A2(g9052B),.A1(g1730B));
AND2_X1 U_g9660B (.ZN(g9660B),.A2(FE_OFN45_g9125B),.A1(g1188B));
AND2_X1 U_g9946B (.ZN(g9946B),.A2(FE_OFN68_g9392B),.A1(g9926B));
AND2_X1 U_g5257B (.ZN(g5257B),.A2(FE_OFN335_g4737B),.A1(g691B));
AND2_X1 U_g4732B (.ZN(g4732B),.A2(FE_OFN300_g4002B),.A1(g391B));
AND2_X1 U_g3108B (.ZN(g3108B),.A2(I6331B),.A1(I6330B));
AND2_X1 U_g4753B (.ZN(g4753B),.A2(FE_OFN307_g4010B),.A1(g481B));
AND2_X1 U_g9903B (.ZN(g9903B),.A2(g9673B),.A1(g9885B));
AND2_X1 U_g10625B (.ZN(g10625B),.A2(FE_OFN369_g4525B),.A1(g10454B));
AND2_X1 U_g5605B (.ZN(g5605B),.A2(g704B),.A1(g4828B));
AND2_X1 U_g6623B (.ZN(g6623B),.A2(FE_OFN97_I8869B),.A1(g55B));
AND2_X1 U_g11228B (.ZN(g11228B),.A2(g11060B),.A1(g466B));
AND2_X1 U_g11011B (.ZN(g11011B),.A2(g10809B),.A1(g1968B));
AND2_X1 U_g6889B (.ZN(g6889B),.A2(FE_OFN213_g6003B),.A1(g1941B));
AND2_X1 U_g8040B (.ZN(g8040B),.A2(FE_OFN305_g5151B),.A1(g7523B));
AND2_X1 U_g7822B (.ZN(g7822B),.A2(FE_OFN209_g6863B),.A1(g1914B));
AND2_X1 U_g8123B (.ZN(g8123B),.A2(g7952B),.A1(g1918B));
AND2_X1 U_g11582B (.ZN(g11582B),.A2(g11539B),.A1(g1311B));
AND2_X1 U_g4316B (.ZN(g4316B),.A2(g3275B),.A1(g1965B));
AND2_X1 U_g10969B (.ZN(g10969B),.A2(g10809B),.A1(g3625B));
AND2_X1 U_g5041B (.ZN(g5041B),.A2(FE_OFN223_g4401B),.A1(g3983B));
AND2_X1 U_g9335B (.ZN(g9335B),.A2(FE_OFN275_g48B),.A1(g8975B));
AND2_X1 U_g9831B (.ZN(g9831B),.A2(FE_OFN34_g9785B),.A1(g9727B));
AND2_X1 U_g4565B (.ZN(g4565B),.A2(g4010B),.A1(g534B));
AND2_X1 U_g9422B (.ZN(g9422B),.A2(FE_OFN50_g9030B),.A1(g1750B));
AND2_X1 U_g8648B (.ZN(g8648B),.A2(g8511B),.A1(g4588B));
AND3_X1 U_g8875B (.ZN(g8875B),.A3(g8858B),.A2(FE_OFN92_g2216B),.A1(g8255B));
AND2_X1 U_g5168B (.ZN(g5168B),.A2(g4679B),.A1(g1512B));
AND2_X1 U_g7895B (.ZN(g7895B),.A2(FE_OFN334_g7045B),.A1(g7503B));
AND2_X1 U_g8655B (.ZN(g8655B),.A2(FE_OFN298_g3015B),.A1(g8267B));
AND2_X1 U_g4914B (.ZN(g4914B),.A2(FE_OFN290_g4880B),.A1(g1062B));
AND2_X1 U_g9947B (.ZN(g9947B),.A2(g9392B),.A1(g9927B));
AND2_X1 U_g5772B (.ZN(g5772B),.A2(FE_OFN321_g5261B),.A1(g1555B));
AND2_X1 U_g6838B (.ZN(g6838B),.A2(FE_OFN180_g5354B),.A1(g192B));
AND2_X1 U_g5531B (.ZN(g5531B),.A2(g4290B),.A1(g1666B));
AND2_X1 U_g6795B (.ZN(g6795B),.A2(g5878B),.A1(g5036B));
AND2_X1 U_g10503B (.ZN(g10503B),.A2(FE_OFN336_g1690B),.A1(g9995B));
AND2_X1 U_g8010B (.ZN(g8010B),.A2(g7438B),.A1(g7738B));
AND2_X1 U_g8410B (.ZN(g8410B),.A2(g8146B),.A1(g713B));
AND2_X1 U_g6231B (.ZN(g6231B),.A2(g5608B),.A1(g818B));
AND2_X1 U_g10581B (.ZN(g10581B),.A2(g9473B),.A1(g10336B));
AND2_X1 U_g10450B (.ZN(g10450B),.A2(FE_OFN235_g2024B),.A1(g10364B));
AND2_X1 U_g2804B (.ZN(g2804B),.A2(g1891B),.A1(g2132B));
AND2_X1 U_g3418B (.ZN(g3418B),.A2(FE_OFN352_g109B),.A1(g2379B));
AND2_X1 U_g9653B (.ZN(g9653B),.A2(FE_OFN45_g9125B),.A1(g1185B));
AND2_X1 U_g6205B (.ZN(g6205B),.A2(FE_OFN306_g5128B),.A1(g1515B));
AND2_X1 U_g10818B (.ZN(g10818B),.A2(FE_OFN204_g3664B),.A1(I16220B));
AND2_X1 U_g8172B (.ZN(g8172B),.A2(FE_OFN89_I11360B),.A1(g37B));
AND2_X1 U_g10496B (.ZN(g10496B),.A2(FE_OFN234_g2024B),.A1(g10429B));
AND2_X1 U_g5074B (.ZN(g5074B),.A2(g4608B),.A1(g1771B));
AND2_X1 U_g9869B (.ZN(g9869B),.A2(g9814B),.A1(g1558B));
AND2_X1 U_g9719B (.ZN(g9719B),.A2(g9490B),.A1(g1543B));
AND2_X1 U_g10741B (.ZN(g10741B),.A2(FE_OFN133_g3015B),.A1(g10635B));
AND2_X1 U_g3381B (.ZN(g3381B),.A2(g2756B),.A1(g940B));
AND2_X1 U_g5863B (.ZN(g5863B),.A2(g622B),.A1(g255B));
AND2_X1 U_g8693B (.ZN(g8693B),.A2(g8509B),.A1(g3738B));
AND2_X1 U_g5480B (.ZN(g5480B),.A2(FE_OFN366_g3521B),.A1(g554B));
AND2_X1 U_g4581B (.ZN(g4581B),.A2(g2047B),.A1(g3766B));
AND2_X1 U_g3685B (.ZN(g3685B),.A2(g2981B),.A1(FE_OFN238_g1781B));
AND2_X1 U_g5569B (.ZN(g5569B),.A2(g2338B),.A1(g4816B));
AND2_X1 U_g8555B (.ZN(g8555B),.A2(FE_OFN189_g7638B),.A1(g8409B));
AND2_X1 U_g3263B (.ZN(g3263B),.A2(g2328B),.A1(g2503B));
AND2_X1 U_g9364B (.ZN(g9364B),.A2(g9223B),.A1(g965B));
AND2_X1 U_g4784B (.ZN(g4784B),.A2(FE_OFN307_g4010B),.A1(g506B));
AND2_X4 U_g9454B (.ZN(g9454B),.A2(FE_OFN275_g48B),.A1(g8994B));
AND4_X1 U_I6331B (.ZN(I6331B),.A4(g2077B),.A3(g2074B),.A2(g2070B),.A1(g2060B));
AND2_X1 U_g11299B (.ZN(g11299B),.A2(g11243B),.A1(g4576B));
AND2_X1 U_g6983B (.ZN(g6983B),.A2(FE_OFN343_I5565B),.A1(g6592B));
AND2_X1 U_g7958B (.ZN(g7958B),.A2(FE_OFN198_g7697B),.A1(g736B));
AND2_X1 U_g4995B (.ZN(g4995B),.A2(FE_OFN153_g4640B),.A1(g1474B));
AND2_X1 U_g4079B (.ZN(g4079B),.A2(g2276B),.A1(FE_OFN237_g1806B));
AND2_X1 U_g2264B (.ZN(g2264B),.A2(g1766B),.A1(FE_OFN247_g1771B));
AND2_X1 U_g2160B (.ZN(g2160B),.A2(g746B),.A1(g745B));
AND2_X1 U_g3257B (.ZN(g3257B),.A2(g2496B),.A1(g378B));
AND2_X1 U_g3101B (.ZN(g3101B),.A2(I6310B),.A1(I6309B));
AND2_X1 U_g5000B (.ZN(g5000B),.A2(FE_OFN153_g4640B),.A1(g1470B));
AND2_X1 U_g3301B (.ZN(g3301B),.A2(g2544B),.A1(g1346B));
AND2_X1 U_g5126B (.ZN(g5126B),.A2(g4671B),.A1(g1104B));
AND4_X1 U_I5084B (.ZN(I5084B),.A4(g1478B),.A3(g1474B),.A2(g1470B),.A1(g1462B));
AND2_X1 U_g9412B (.ZN(g9412B),.A2(g9052B),.A1(g1727B));
AND2_X1 U_g9389B (.ZN(g9389B),.A2(FE_OFN47_g9151B),.A1(g1330B));
AND2_X1 U_g2379B (.ZN(g2379B),.A2(g743B),.A1(g744B));
AND2_X1 U_g10706B (.ZN(g10706B),.A2(FE_OFN345_g3015B),.A1(g10567B));
AND3_X1 U_I16145B (.ZN(I16145B),.A3(g10446B),.A2(g10447B),.A1(g10366B));
AND2_X1 U_g10597B (.ZN(g10597B),.A2(FE_OFN369_g4525B),.A1(g10533B));
AND3_X1 U_g8965B (.ZN(g8965B),.A3(g8849B),.A2(FE_OFN281_g2216B),.A1(g8110B));
AND2_X1 U_g5608B (.ZN(g5608B),.A2(g4831B),.A1(g814B));
AND2_X1 U_g5220B (.ZN(g5220B),.A2(g4776B),.A1(g1083B));
AND2_X1 U_g10624B (.ZN(g10624B),.A2(FE_OFN370_g4525B),.A1(g10494B));
AND2_X1 U_g10300B (.ZN(g10300B),.A2(g10019B),.A1(FE_OFN76_g8700B));
AND2_X1 U_g5023B (.ZN(g5023B),.A2(FE_OFN288_g4263B),.A1(g1071B));
AND2_X1 U_g4432B (.ZN(g4432B),.A2(g1975B),.A1(g3723B));
AND2_X1 U_g4053B (.ZN(g4053B),.A2(FE_OFN224_g2276B),.A1(FE_OFN253_g1786B));
AND2_X1 U_g8050B (.ZN(g8050B),.A2(FE_OFN177_g5919B),.A1(g7596B));
AND2_X1 U_g5588B (.ZN(g5588B),.A2(FE_OFN367_g3521B),.A1(g1639B));
AND3_X1 U_g6679B (.ZN(g6679B),.A3(g109B),.A2(g6074B),.A1(FE_OFN184_I7048B));
AND2_X1 U_g9963B (.ZN(g9963B),.A2(FE_OFN280_g9536B),.A1(g9953B));
AND2_X1 U_g3772B (.ZN(g3772B),.A2(g3089B),.A1(g2542B));
AND2_X1 U_g5051B (.ZN(g5051B),.A2(g2506B),.A1(g4432B));
AND2_X1 U_g6831B (.ZN(g6831B),.A2(FE_OFN179_g5354B),.A1(g207B));
AND2_X1 U_g2981B (.ZN(g2981B),.A2(g2264B),.A1(FE_OFN236_g1776B));
AND2_X1 U_g8724B (.ZN(g8724B),.A2(g7910B),.A1(g8214B));
AND2_X1 U_g4157B (.ZN(g4157B),.A2(g3060B),.A1(FE_OFN239_g1796B));
AND2_X1 U_g9707B (.ZN(g9707B),.A2(g9474B),.A1(g1583B));
AND3_X1 U_g8878B (.ZN(g8878B),.A3(FE_OFN73_g8858B),.A2(FE_OFN93_g2216B),.A1(g8099B));
AND2_X1 U_g2132B (.ZN(g2132B),.A2(g1882B),.A1(g1872B));
AND2_X1 U_g10763B (.ZN(g10763B),.A2(FE_OFN345_g3015B),.A1(g10639B));
AND3_X1 U_g8289B (.ZN(g8289B),.A3(g2216B),.A2(g8109B),.A1(g6777B));
AND2_X1 U_g7898B (.ZN(g7898B),.A2(g7045B),.A1(g7511B));
AND2_X1 U_g11271B (.ZN(g11271B),.A2(g11203B),.A1(g4753B));
AND2_X1 U_g11461B (.ZN(g11461B),.A2(FE_OFN100_g4421B),.A1(g11225B));
AND2_X1 U_g5732B (.ZN(g5732B),.A2(FE_OFN353_g5117B),.A1(g1604B));
AND2_X1 U_g11145B (.ZN(g11145B),.A2(FE_OFN278_g10927B),.A1(g315B));
AND2_X1 U_g11031B (.ZN(g11031B),.A2(FE_OFN14_g10702B),.A1(g411B));
AND2_X1 U_g9865B (.ZN(g9865B),.A2(g9773B),.A1(g1607B));
AND2_X1 U_g5944B (.ZN(g5944B),.A2(g5233B),.A1(g1796B));
AND2_X1 U_g9715B (.ZN(g9715B),.A2(FE_OFN70_g9490B),.A1(g1531B));
AND2_X1 U_g9604B (.ZN(g9604B),.A2(FE_OFN51_g9111B),.A1(g1194B));
AND2_X1 U_g8799B (.ZN(g8799B),.A2(FE_OFN331_g8696B),.A1(g8647B));
AND2_X1 U_g11198B (.ZN(g11198B),.A2(FE_OFN15_g10702B),.A1(g4778B));
AND2_X1 U_g6873B (.ZN(g6873B),.A2(g6557B),.A1(g3263B));
AND2_X1 U_g6632B (.ZN(g6632B),.A2(FE_OFN283_I8869B),.A1(g61B));
AND2_X1 U_g6095B (.ZN(g6095B),.A2(FE_OFN273_g85B),.A1(g1062B));
AND2_X1 U_g3863B (.ZN(g3863B),.A2(g1696B),.A1(g1703B));
AND2_X1 U_g9833B (.ZN(g9833B),.A2(FE_OFN34_g9785B),.A1(g9729B));
AND2_X1 U_g6653B (.ZN(g6653B),.A2(I8869B),.A1(g70B));
AND2_X1 U_g6102B (.ZN(g6102B),.A2(FE_OFN273_g85B),.A1(g1038B));
AND2_X1 U_g7819B (.ZN(g7819B),.A2(FE_OFN206_g6863B),.A1(g1887B));
AND2_X1 U_g11393B (.ZN(g11393B),.A2(g7914B),.A1(g11280B));
AND2_X1 U_g2511B (.ZN(g2511B),.A2(g456B),.A1(FE_OFN254_g461B));
AND2_X1 U_g7088B (.ZN(g7088B),.A2(g6432B),.A1(g2331B));
AND2_X1 U_g9584B (.ZN(g9584B),.A2(FE_OFN53_g9173B),.A1(g1341B));
AND2_X1 U_g9896B (.ZN(g9896B),.A2(FE_OFN60_g9624B),.A1(g9696B));
AND3_X1 U_g8209B (.ZN(g8209B),.A3(g7622B),.A2(g3068B),.A1(g4094B));
AND2_X1 U_g6752B (.ZN(g6752B),.A2(g2343B),.A1(g6187B));
AND2_X1 U_g4778B (.ZN(g4778B),.A2(g4002B),.A1(g421B));
AND2_X1 U_g11161B (.ZN(g11161B),.A2(g10937B),.A1(g1969B));
AND2_X1 U_g9268B (.ZN(g9268B),.A2(g8947B),.A1(g6109B));
AND2_X1 U_g5681B (.ZN(g5681B),.A2(FE_OFN365_g5361B),.A1(g135B));
AND2_X1 U_g7951B (.ZN(g7951B),.A2(g7505B),.A1(g73B));
AND2_X1 U_g9419B (.ZN(g9419B),.A2(FE_OFN50_g9030B),.A1(g1744B));
AND2_X1 U_g10268B (.ZN(g10268B),.A2(FE_OFN267_g109B),.A1(I15287B));
AND2_X1 U_g5533B (.ZN(g5533B),.A2(g4292B),.A1(g1724B));
AND2_X4 U_g9052B (.ZN(g9052B),.A2(FE_OFN276_g48B),.A1(g8936B));
AND2_X1 U_g6786B (.ZN(g6786B),.A2(g5919B),.A1(g178B));
AND2_X1 U_g10670B (.ZN(g10670B),.A2(g9097B),.A1(g10396B));
AND2_X1 U_g11087B (.ZN(g11087B),.A2(FE_OFN4_g10950B),.A1(g829B));
AND2_X1 U_g4949B (.ZN(g4949B),.A2(g4449B),.A1(I5815B));
AND2_X1 U_g6364B (.ZN(g6364B),.A2(FE_OFN346_g4381B),.A1(g5851B));
AND2_X1 U_g7825B (.ZN(g7825B),.A2(FE_OFN206_g6863B),.A1(g1941B));
AND2_X1 U_g4998B (.ZN(g4998B),.A2(FE_OFN303_g4678B),.A1(g1304B));
AND2_X1 U_g10667B (.ZN(g10667B),.A2(g9424B),.A1(g10405B));
AND2_X1 U_g7136B (.ZN(g7136B),.A2(g6718B),.A1(g5190B));
AND2_X1 U_g6532B (.ZN(g6532B),.A2(FE_OFN282_g6165B),.A1(g339B));
AND2_X1 U_g9385B (.ZN(g9385B),.A2(FE_OFN48_g9151B),.A1(g1324B));
AND4_X1 U_I5690B (.ZN(I5690B),.A4(g1448B),.A3(g1444B),.A2(g1440B),.A1(g1436B));
AND2_X1 U_g4484B (.ZN(g4484B),.A2(FE_OFN302_g3913B),.A1(g1137B));
AND2_X1 U_g9897B (.ZN(g9897B),.A2(FE_OFN60_g9624B),.A1(g9699B));
AND2_X1 U_g9425B (.ZN(g9425B),.A2(FE_OFN49_g9030B),.A1(g1753B));
AND2_X1 U_g3383B (.ZN(g3383B),.A2(FE_OFN324_g18B),.A1(g186B));
AND2_X1 U_g5601B (.ZN(g5601B),.A2(g4880B),.A1(g1035B));
AND2_X1 U_g7943B (.ZN(g7943B),.A2(g7467B),.A1(g64B));
AND2_X1 U_g11171B (.ZN(g11171B),.A2(FE_OFN21_g10702B),.A1(g481B));
AND2_X1 U_g3423B (.ZN(g3423B),.A2(I6631B),.A1(I6630B));
AND2_X1 U_g7230B (.ZN(g7230B),.A2(g6447B),.A1(g6064B));
AND2_X1 U_g4952B (.ZN(g4952B),.A2(FE_OFN299_g4457B),.A1(g1648B));
AND2_X1 U_g6787B (.ZN(g6787B),.A2(FE_OFN319_g5361B),.A1(g266B));
AND3_X1 U_g8968B (.ZN(g8968B),.A3(g8849B),.A2(FE_OFN281_g2216B),.A1(g8089B));
AND2_X1 U_g10306B (.ZN(g10306B),.A2(g9082B),.A1(g10007B));
AND2_X1 U_g9331B (.ZN(g9331B),.A2(FE_OFN275_g48B),.A1(g8972B));
AND2_X1 U_g11459B (.ZN(g11459B),.A2(FE_OFN100_g4421B),.A1(g11221B));
AND2_X1 U_g4561B (.ZN(g4561B),.A2(g4010B),.A1(g538B));
AND2_X1 U_g11425B (.ZN(g11425B),.A2(g10629B),.A1(I16982B));
AND2_X1 U_g11458B (.ZN(g11458B),.A2(FE_OFN99_g4421B),.A1(g11219B));
AND2_X1 U_g5739B (.ZN(g5739B),.A2(FE_OFN315_g5117B),.A1(g1607B));
AND2_X1 U_g7496B (.ZN(g7496B),.A2(g64B),.A1(FE_OFN83_g2176B));
AND2_X1 U_g4986B (.ZN(g4986B),.A2(FE_OFN146_g4682B),.A1(g1411B));
AND2_X1 U_g11010B (.ZN(g11010B),.A2(FE_OFN18_g10702B),.A1(g5187B));
AND2_X1 U_g3999B (.ZN(g3999B),.A2(g2777B),.A1(g1741B));
AND2_X1 U_g8175B (.ZN(g8175B),.A2(FE_OFN89_I11360B),.A1(g39B));
AND2_X1 U_g8722B (.ZN(g8722B),.A2(g7908B),.A1(g8210B));
AND2_X1 U_g4764B (.ZN(g4764B),.A2(FE_OFN300_g4002B),.A1(g411B));
AND2_X1 U_g7137B (.ZN(g7137B),.A2(g6354B),.A1(g5590B));
AND2_X1 U_g7891B (.ZN(g7891B),.A2(FE_OFN334_g7045B),.A1(g7471B));
AND2_X1 U_g8651B (.ZN(g8651B),.A2(FE_OFN348_g3015B),.A1(g8261B));
AND2_X1 U_g5479B (.ZN(g5479B),.A2(g4243B),.A1(g1845B));
AND2_X1 U_g11599B (.ZN(g11599B),.A2(g11575B),.A1(g1341B));
AND2_X1 U_g6684B (.ZN(g6684B),.A2(g5836B),.A1(g91B));
AND2_X1 U_g6745B (.ZN(g6745B),.A2(FE_OFN218_g5557B),.A1(g5605B));
AND2_X1 U_g6639B (.ZN(g6639B),.A2(FE_OFN282_g6165B),.A1(g357B));
AND2_X1 U_g10937B (.ZN(g10937B),.A2(FE_OFN13_g10702B),.A1(g4822B));
AND2_X1 U_g3696B (.ZN(g3696B),.A2(FE_OFN364_g3015B),.A1(g1713B));
AND2_X1 U_g4503B (.ZN(g4503B),.A2(g3943B),.A1(g654B));
AND2_X1 U_g6791B (.ZN(g6791B),.A2(FE_OFN319_g5361B),.A1(g269B));
AND2_X1 U_g5190B (.ZN(g5190B),.A2(g4678B),.A1(g1245B));
AND2_X1 U_g5390B (.ZN(g5390B),.A2(g4671B),.A1(g1101B));
AND2_X1 U_g8384B (.ZN(g8384B),.A2(FE_OFN325_g18B),.A1(g8180B));
AND2_X1 U_g4224B (.ZN(g4224B),.A2(FE_OFN132_g3015B),.A1(g1092B));
AND2_X1 U_g5501B (.ZN(g5501B),.A2(g4273B),.A1(g1672B));
AND2_X4 U_g9173B (.ZN(g9173B),.A2(FE_OFN276_g48B),.A1(g8968B));
AND2_X1 U_g6759B (.ZN(g6759B),.A2(g5919B),.A1(g148B));
AND2_X1 U_g8838B (.ZN(g8838B),.A2(FE_OFN328_g8709B),.A1(g8602B));
AND2_X1 U_g8024B (.ZN(g8024B),.A2(FE_OFN322_g4449B),.A1(g6577B));
AND2_X1 U_g10666B (.ZN(g10666B),.A2(g9424B),.A1(g10402B));
AND2_X1 U_g11158B (.ZN(g11158B),.A2(FE_OFN278_g10927B),.A1(g309B));
AND2_X1 U_g9602B (.ZN(g9602B),.A2(g9010B),.A1(g932B));
AND2_X1 U_g5704B (.ZN(g5704B),.A2(FE_OFN164_g5361B),.A1(g143B));
AND2_X1 U_g4617B (.ZN(g4617B),.A2(g3879B),.A1(g3275B));
AND2_X2 U_g11561B (.ZN(g11561B),.A2(FE_OFN364_g3015B),.A1(g11492B));
AND2_X1 U_g9868B (.ZN(g9868B),.A2(g9814B),.A1(g1555B));
AND2_X1 U_g11295B (.ZN(g11295B),.A2(g11239B),.A1(g4554B));
AND2_X1 U_g11144B (.ZN(g11144B),.A2(FE_OFN10_g10702B),.A1(g305B));
AND2_X1 U_g9718B (.ZN(g9718B),.A2(FE_OFN70_g9490B),.A1(g1540B));
AND2_X1 U_g3434B (.ZN(g3434B),.A2(g2355B),.A1(g237B));
AND2_X1 U_g4987B (.ZN(g4987B),.A2(FE_OFN147_g4682B),.A1(g1440B));
AND2_X1 U_g4771B (.ZN(g4771B),.A2(FE_OFN307_g4010B),.A1(g496B));
AND2_X1 U_g5250B (.ZN(g5250B),.A2(g4678B),.A1(g1270B));
AND2_X1 U_g6098B (.ZN(g6098B),.A2(FE_OFN273_g85B),.A1(g1065B));
AND2_X1 U_g9582B (.ZN(g9582B),.A2(FE_OFN53_g9173B),.A1(g2725B));
AND2_X1 U_g6833B (.ZN(g6833B),.A2(FE_OFN178_g5354B),.A1(g186B));
AND2_X1 U_g3533B (.ZN(g3533B),.A2(g2892B),.A1(g1981B));
AND2_X1 U_g4892B (.ZN(g4892B),.A2(g4739B),.A1(g632B));
AND2_X1 U_g8104B (.ZN(g8104B),.A2(g7852B),.A1(g5493B));
AND2_X1 U_g9415B (.ZN(g9415B),.A2(FE_OFN54_g9052B),.A1(g1733B));
AND2_X1 U_g8499B (.ZN(g8499B),.A2(g4737B),.A1(g8377B));
AND2_X1 U_g9664B (.ZN(g9664B),.A2(FE_OFN46_g9125B),.A1(g1191B));
AND2_X1 U_g9721B (.ZN(g9721B),.A2(FE_OFN359_g18B),.A1(g9413B));
AND2_X1 U_g6162B (.ZN(g6162B),.A2(g5200B),.A1(g3584B));
AND2_X1 U_g4991B (.ZN(g4991B),.A2(FE_OFN154_g4640B),.A1(g1508B));
AND2_X1 U_g6362B (.ZN(g6362B),.A2(FE_OFN346_g4381B),.A1(g5846B));
AND4_X1 U_I6631B (.ZN(I6631B),.A4(FE_OFN237_g1806B),.A3(FE_OFN251_g1801B),.A2(FE_OFN239_g1796B),.A1(FE_OFN252_g1791B));
AND2_X1 U_g10685B (.ZN(g10685B),.A2(FE_OFN136_g3863B),.A1(g10383B));
AND2_X1 U_g4340B (.ZN(g4340B),.A2(FE_OFN351_g3913B),.A1(g1153B));
AND2_X1 U_g11023B (.ZN(g11023B),.A2(g10702B),.A1(g440B));
AND2_X1 U_g8044B (.ZN(g8044B),.A2(FE_OFN177_g5919B),.A1(g7598B));
AND2_X1 U_g11224B (.ZN(g11224B),.A2(g11157B),.A1(g968B));
AND2_X1 U_g11571B (.ZN(g11571B),.A2(g11561B),.A1(g2018B));
AND2_X1 U_g4959B (.ZN(g4959B),.A2(FE_OFN147_g4682B),.A1(g1520B));
AND2_X1 U_g10334B (.ZN(g10334B),.A2(FE_OFN267_g109B),.A1(I15365B));
AND2_X1 U_g5626B (.ZN(g5626B),.A2(FE_OFN367_g3521B),.A1(g1633B));
AND2_X1 U_g9940B (.ZN(g9940B),.A2(FE_OFN67_g9367B),.A1(g9920B));
AND2_X1 U_g4876B (.ZN(g4876B),.A2(FE_OFN132_g3015B),.A1(g1086B));
AND2_X1 U_g6728B (.ZN(g6728B),.A2(FE_OFN310_g4336B),.A1(g4482B));
AND2_X1 U_g6730B (.ZN(g6730B),.A2(g5013B),.A1(g1872B));
AND2_X1 U_g9689B (.ZN(g9689B),.A2(FE_OFN59_g9432B),.A1(g263B));
AND2_X1 U_g10762B (.ZN(g10762B),.A2(FE_OFN131_g3015B),.A1(g10635B));
AND2_X1 U_g6070B (.ZN(g6070B),.A2(FE_OFN273_g85B),.A1(g1050B));
AND2_X1 U_g9428B (.ZN(g9428B),.A2(FE_OFN50_g9030B),.A1(g1756B));
AND2_X4 U_g9030B (.ZN(g9030B),.A2(FE_OFN276_g48B),.A1(g8935B));
AND2_X1 U_g9430B (.ZN(g9430B),.A2(FE_OFN49_g9030B),.A1(g1759B));
AND2_X1 U_g8927B (.ZN(g8927B),.A2(g8642B),.A1(g2216B));
AND2_X1 U_g7068B (.ZN(g7068B),.A2(g6586B),.A1(g5024B));
AND2_X1 U_g8014B (.ZN(g8014B),.A2(g7438B),.A1(g7740B));
AND2_X1 U_g11392B (.ZN(g11392B),.A2(g7914B),.A1(g11278B));
AND2_X1 U_g5782B (.ZN(g5782B),.A2(g5222B),.A1(g1558B));
AND2_X1 U_g4824B (.ZN(g4824B),.A2(g4099B),.A1(g774B));
AND2_X1 U_g6331B (.ZN(g6331B),.A2(FE_OFN180_g5354B),.A1(g201B));
AND2_X1 U_g4236B (.ZN(g4236B),.A2(FE_OFN132_g3015B),.A1(g1098B));
AND2_X1 U_g11559B (.ZN(g11559B),.A2(FE_OFN27_g11519B),.A1(FE_OFN251_g1801B));
AND2_X1 U_g9609B (.ZN(g9609B),.A2(FE_OFN42_g9205B),.A1(g907B));
AND2_X1 U_g11558B (.ZN(g11558B),.A2(FE_OFN27_g11519B),.A1(FE_OFN239_g1796B));
AND2_X1 U_g6087B (.ZN(g6087B),.A2(FE_OFN271_g85B),.A1(g1056B));
AND2_X1 U_g5526B (.ZN(g5526B),.A2(g4294B),.A1(g1950B));
AND2_X1 U_g10751B (.ZN(g10751B),.A2(FE_OFN133_g3015B),.A1(g10646B));
AND2_X1 U_g10772B (.ZN(g10772B),.A2(FE_OFN345_g3015B),.A1(g10655B));
AND2_X1 U_g8135B (.ZN(g8135B),.A2(g7883B),.A1(g1945B));
AND2_X1 U_g11544B (.ZN(g11544B),.A2(g10584B),.A1(g11515B));
AND2_X1 U_g5084B (.ZN(g5084B),.A2(FE_OFN299_g4457B),.A1(g1776B));
AND2_X1 U_g8382B (.ZN(g8382B),.A2(FE_OFN196_g7697B),.A1(g5248B));
AND2_X1 U_g10230B (.ZN(g10230B),.A2(g9968B),.A1(g8700B));
AND2_X1 U_g5484B (.ZN(g5484B),.A2(FE_OFN333_g4294B),.A1(g1896B));
AND2_X1 U_g7241B (.ZN(g7241B),.A2(g5557B),.A1(g6772B));
AND2_X1 U_g3942B (.ZN(g3942B),.A2(FE_OFN260_g18B),.A1(g219B));
AND2_X1 U_g10638B (.ZN(g10638B),.A2(g3829B),.A1(g10383B));
AND2_X1 U_g4064B (.ZN(g4064B),.A2(g2774B),.A1(g1759B));
AND2_X1 U_g9365B (.ZN(g9365B),.A2(FE_OFN48_g9151B),.A1(g1321B));
AND2_X1 U_g9861B (.ZN(g9861B),.A2(g9579B),.A1(g9738B));
AND2_X1 U_g11255B (.ZN(g11255B),.A2(g11060B),.A1(g456B));
AND2_X1 U_g11189B (.ZN(g11189B),.A2(FE_OFN15_g10702B),.A1(g4736B));
AND2_X1 U_g10510B (.ZN(g10510B),.A2(FE_OFN336_g1690B),.A1(g10019B));
AND3_X1 U_g8947B (.ZN(g8947B),.A3(g8828B),.A2(FE_OFN92_g2216B),.A1(g8056B));
AND2_X1 U_g2917B (.ZN(g2917B),.A2(g1657B),.A1(g2424B));
AND2_X2 U_g5919B (.ZN(g5919B),.A2(FE_OFN269_g109B),.A1(I7048B));
AND2_X1 U_g11188B (.ZN(g11188B),.A2(FE_OFN15_g10702B),.A1(g4732B));
AND2_X1 U_g9846B (.ZN(g9846B),.A2(g9764B),.A1(g287B));
AND2_X1 U_g7818B (.ZN(g7818B),.A2(FE_OFN206_g6863B),.A1(g1878B));
AND2_X1 U_g11460B (.ZN(g11460B),.A2(FE_OFN99_g4421B),.A1(g11223B));
AND2_X1 U_g5276B (.ZN(g5276B),.A2(FE_OFN335_g4737B),.A1(g736B));
AND2_X1 U_g11030B (.ZN(g11030B),.A2(FE_OFN17_g10702B),.A1(g406B));
AND2_X1 U_g11093B (.ZN(g11093B),.A2(FE_OFN4_g10950B),.A1(g841B));
AND2_X1 U_g7893B (.ZN(g7893B),.A2(FE_OFN334_g7045B),.A1(g7478B));
AND2_X1 U_g8653B (.ZN(g8653B),.A2(FE_OFN348_g3015B),.A1(g8265B));
AND2_X1 U_g10442B (.ZN(g10442B),.A2(FE_OFN245_g1690B),.A1(g9968B));
AND2_X1 U_g6535B (.ZN(g6535B),.A2(g6165B),.A1(g345B));
AND2_X1 U_g8102B (.ZN(g8102B),.A2(g7852B),.A1(g5485B));
AND4_X1 U_I5085B (.ZN(I5085B),.A4(g1508B),.A3(g1504B),.A2(g1494B),.A1(g1490B));
AND2_X1 U_g5004B (.ZN(g5004B),.A2(FE_OFN303_g4678B),.A1(g1296B));
AND2_X1 U_g3912B (.ZN(g3912B),.A2(FE_OFN359_g18B),.A1(g207B));
AND2_X1 U_g7186B (.ZN(g7186B),.A2(g6403B),.A1(g2503B));
AND2_X1 U_g4489B (.ZN(g4489B),.A2(FE_OFN103_g3586B),.A1(g348B));
AND2_X1 U_g9662B (.ZN(g9662B),.A2(g9292B),.A1(g123B));
AND2_X1 U_g9418B (.ZN(g9418B),.A2(FE_OFN56_g9052B),.A1(g1741B));
AND2_X1 U_g11218B (.ZN(g11218B),.A2(FE_OFN279_g11157B),.A1(g959B));
AND2_X1 U_g4471B (.ZN(g4471B),.A2(FE_OFN302_g3913B),.A1(g1121B));
AND2_X1 U_g10746B (.ZN(g10746B),.A2(FE_OFN364_g3015B),.A1(g10643B));
AND2_X1 U_g7125B (.ZN(g7125B),.A2(g5763B),.A1(g1212B));
AND2_X1 U_g7821B (.ZN(g7821B),.A2(FE_OFN209_g6863B),.A1(g1905B));
AND2_X1 U_g6246B (.ZN(g6246B),.A2(FE_OFN164_g5361B),.A1(g178B));
AND2_X1 U_g9256B (.ZN(g9256B),.A2(g8963B),.A1(g6109B));
AND2_X1 U_g8042B (.ZN(g8042B),.A2(FE_OFN305_g5151B),.A1(g7533B));
AND2_X1 U_g10237B (.ZN(g10237B),.A2(g9082B),.A1(g9968B));
AND2_X1 U_g7939B (.ZN(g7939B),.A2(g7460B),.A1(g61B));
AND2_X1 U_g8786B (.ZN(g8786B),.A2(FE_OFN331_g8696B),.A1(g8638B));
AND2_X1 U_g10684B (.ZN(g10684B),.A2(FE_OFN136_g3863B),.A1(g10382B));
AND2_X1 U_g11455B (.ZN(g11455B),.A2(FE_OFN99_g4421B),.A1(g11233B));
AND2_X1 U_g8364B (.ZN(g8364B),.A2(g8146B),.A1(g658B));
AND3_X1 U_g2990B (.ZN(g2990B),.A3(g1814B),.A2(g2557B),.A1(g2061B));
AND2_X1 U_g9847B (.ZN(g9847B),.A2(FE_OFN57_g9432B),.A1(g290B));
AND2_X1 U_g8054B (.ZN(g8054B),.A2(FE_OFN177_g5919B),.A1(g7584B));
AND2_X1 U_g5617B (.ZN(g5617B),.A2(FE_OFN290_g4880B),.A1(g1050B));
AND2_X1 U_g6502B (.ZN(g6502B),.A2(FE_OFN363_I5565B),.A1(g5981B));
AND2_X1 U_g5789B (.ZN(g5789B),.A2(FE_OFN321_g5261B),.A1(g1561B));
AND2_X1 U_g4009B (.ZN(g4009B),.A2(g2774B),.A1(g1747B));
AND2_X1 U_g11277B (.ZN(g11277B),.A2(g11199B),.A1(g4779B));
AND2_X1 U_g6940B (.ZN(g6940B),.A2(g1945B),.A1(g6472B));
AND2_X1 U_g7061B (.ZN(g7061B),.A2(g6760B),.A1(g790B));
AND2_X1 U_g11595B (.ZN(g11595B),.A2(g11575B),.A1(g1336B));
AND2_X1 U_g5771B (.ZN(g5771B),.A2(FE_OFN321_g5261B),.A1(g1534B));
AND2_X1 U_g8553B (.ZN(g8553B),.A2(FE_OFN330_g7638B),.A1(g8405B));
AND2_X1 U_g4836B (.ZN(g4836B),.A2(g3943B),.A1(g643B));
AND2_X1 U_g5547B (.ZN(g5547B),.A2(g4292B),.A1(g1733B));
AND2_X1 U_g6216B (.ZN(g6216B),.A2(FE_OFN306_g5128B),.A1(g1407B));
AND2_X1 U_g4967B (.ZN(g4967B),.A2(FE_OFN146_g4682B),.A1(g1515B));
AND2_X1 U_g6671B (.ZN(g6671B),.A2(FE_OFN282_g6165B),.A1(g342B));
AND2_X1 U_g7200B (.ZN(g7200B),.A2(g6447B),.A1(g3098B));
AND2_X1 U_g3661B (.ZN(g3661B),.A2(g3257B),.A1(g382B));
AND2_X1 U_g7046B (.ZN(g7046B),.A2(g6702B),.A1(g4998B));
AND2_X1 U_g4229B (.ZN(g4229B),.A2(g4673B),.A1(g999B));
AND2_X1 U_g8389B (.ZN(g8389B),.A2(g8220B),.A1(g5263B));
AND2_X1 U_g6430B (.ZN(g6430B),.A2(FE_OFN217_g5013B),.A1(g5044B));
AND2_X1 U_g4993B (.ZN(g4993B),.A2(FE_OFN147_g4682B),.A1(g1448B));
AND2_X1 U_g6247B (.ZN(g6247B),.A2(FE_OFN365_g5361B),.A1(g127B));
AND2_X1 U_g9257B (.ZN(g9257B),.A2(g8964B),.A1(g6109B));
AND2_X1 U_g11170B (.ZN(g11170B),.A2(FE_OFN8_g10702B),.A1(g525B));
AND2_X1 U_g7145B (.ZN(g7145B),.A2(g6718B),.A1(g5250B));
AND2_X1 U_g5738B (.ZN(g5738B),.A2(FE_OFN353_g5117B),.A1(g1586B));
AND2_X1 U_g6826B (.ZN(g6826B),.A2(g5354B),.A1(g225B));
AND2_X1 U_g7191B (.ZN(g7191B),.A2(FE_OFN310_g4336B),.A1(g5219B));
AND2_X1 U_g3998B (.ZN(g3998B),.A2(g2276B),.A1(g2677B));
AND2_X1 U_g6741B (.ZN(g6741B),.A2(FE_OFN219_g5557B),.A1(g3284B));
AND2_X1 U_g5478B (.ZN(g5478B),.A2(FE_OFN333_g4294B),.A1(g1905B));
AND2_X1 U_g11167B (.ZN(g11167B),.A2(FE_OFN8_g10702B),.A1(g538B));
AND2_X1 U_g11194B (.ZN(g11194B),.A2(g10927B),.A1(g4764B));
AND2_X1 U_g11589B (.ZN(g11589B),.A2(g11539B),.A1(g1333B));
AND2_X1 U_g6638B (.ZN(g6638B),.A2(FE_OFN283_I8869B),.A1(g64B));
AND2_X2 U_g4921B (.ZN(g4921B),.A2(g4431B),.A1(g627B));
AND2_X1 U_g7536B (.ZN(g7536B),.A2(g76B),.A1(FE_OFN83_g2176B));
AND2_X1 U_g9585B (.ZN(g9585B),.A2(g8995B),.A1(g889B));
AND2_X1 U_g2957B (.ZN(g2957B),.A2(g1663B),.A1(g2424B));
AND2_X1 U_g11588B (.ZN(g11588B),.A2(g11547B),.A1(g1330B));
AND2_X1 U_g5690B (.ZN(g5690B),.A2(FE_OFN353_g5117B),.A1(g1567B));
AND2_X1 U_g6883B (.ZN(g6883B),.A2(FE_OFN213_g6003B),.A1(g1923B));
AND2_X1 U_g4837B (.ZN(g4837B),.A2(FE_OFN297_g3015B),.A1(g1068B));
AND3_X1 U_g8963B (.ZN(g8963B),.A3(g8849B),.A2(FE_OFN92_g2216B),.A1(g8056B));
AND2_X1 U_g8791B (.ZN(g8791B),.A2(FE_OFN331_g8696B),.A1(g8641B));
AND2_X1 U_g6217B (.ZN(g6217B),.A2(FE_OFN291_g4880B),.A1(g563B));
AND4_X1 U_I6316B (.ZN(I6316B),.A4(g2395B),.A3(g2381B),.A2(g2087B),.A1(g2082B));
AND2_X1 U_g11022B (.ZN(g11022B),.A2(g10702B),.A1(g444B));
AND2_X1 U_g5915B (.ZN(g5915B),.A2(g4977B),.A1(g4168B));
AND2_X1 U_g4788B (.ZN(g4788B),.A2(FE_OFN307_g4010B),.A1(g511B));
AND2_X1 U_g5110B (.ZN(g5110B),.A2(FE_OFN299_g4457B),.A1(FE_OFN237_g1806B));
AND2_X1 U_g11254B (.ZN(g11254B),.A2(g11083B),.A1(g986B));
AND2_X1 U_g6827B (.ZN(g6827B),.A2(FE_OFN178_g5354B),.A1(g219B));
AND3_X1 U_g8957B (.ZN(g8957B),.A3(g8828B),.A2(FE_OFN281_g2216B),.A1(g8081B));
AND2_X1 U_g6333B (.ZN(g6333B),.A2(FE_OFN180_g5354B),.A1(g197B));
AND2_X1 U_g8049B (.ZN(g8049B),.A2(FE_OFN177_g5919B),.A1(g7567B));
AND2_X1 U_g4392B (.ZN(g4392B),.A2(FE_OFN137_g3829B),.A1(g3273B));
AND2_X1 U_g9856B (.ZN(g9856B),.A2(g9773B),.A1(g1592B));
AND2_X1 U_g9411B (.ZN(g9411B),.A2(g9052B),.A1(g1724B));
AND2_X1 U_g5002B (.ZN(g5002B),.A2(FE_OFN154_g4640B),.A1(g1494B));
AND2_X1 U_g11101B (.ZN(g11101B),.A2(FE_OFN4_g10950B),.A1(g857B));
AND2_X1 U_g11177B (.ZN(g11177B),.A2(FE_OFN20_g10702B),.A1(g511B));
AND2_X1 U_g11560B (.ZN(g11560B),.A2(FE_OFN27_g11519B),.A1(g1806B));
AND2_X1 U_g8098B (.ZN(g8098B),.A2(g7852B),.A1(g5478B));
AND2_X1 U_g3970B (.ZN(g3970B),.A2(FE_OFN260_g18B),.A1(g225B));
AND2_X1 U_g4941B (.ZN(g4941B),.A2(FE_OFN290_g4880B),.A1(g1038B));
AND2_X1 U_g10453B (.ZN(g10453B),.A2(FE_OFN234_g2024B),.A1(g10437B));
AND2_X1 U_g5877B (.ZN(g5877B),.A2(g639B),.A1(g4921B));
AND2_X1 U_g6662B (.ZN(g6662B),.A2(FE_OFN282_g6165B),.A1(g366B));
AND2_X1 U_g7935B (.ZN(g7935B),.A2(g7454B),.A1(g58B));
AND2_X1 U_g6067B (.ZN(g6067B),.A2(g85B),.A1(g1047B));
AND4_X1 U_I6317B (.ZN(I6317B),.A4(g2438B),.A3(g2434B),.A2(g2420B),.A1(g2406B));
AND2_X1 U_g9863B (.ZN(g9863B),.A2(FE_OFN56_g9052B),.A1(g9740B));
AND4_X1 U_I5886B (.ZN(I5886B),.A4(g2254B),.A3(g2249B),.A2(g170B),.A1(g174B));
AND2_X1 U_g6994B (.ZN(g6994B),.A2(FE_OFN141_g3829B),.A1(g6758B));
AND2_X1 U_g9713B (.ZN(g9713B),.A2(FE_OFN63_g9474B),.A1(g1589B));
AND2_X1 U_g4431B (.ZN(g4431B),.A2(g3533B),.A1(g2268B));
AND2_X1 U_g4252B (.ZN(g4252B),.A2(FE_OFN347_g3914B),.A1(g1007B));
AND2_X1 U_g11166B (.ZN(g11166B),.A2(FE_OFN9_g10702B),.A1(g542B));
AND2_X1 U_g7130B (.ZN(g7130B),.A2(g6697B),.A1(g5150B));
AND2_X1 U_g11009B (.ZN(g11009B),.A2(FE_OFN18_g10702B),.A1(g5179B));
AND2_X1 U_g7542B (.ZN(g7542B),.A2(g79B),.A1(FE_OFN85_g2176B));
AND2_X1 U_g8019B (.ZN(g8019B),.A2(FE_OFN310_g4336B),.A1(g6573B));
AND2_X1 U_g11008B (.ZN(g11008B),.A2(FE_OFN18_g10702B),.A1(g5171B));
AND2_X1 U_g3516B (.ZN(g3516B),.A2(FE_OFN298_g3015B),.A1(g1209B));
AND2_X1 U_g8052B (.ZN(g8052B),.A2(FE_OFN305_g5151B),.A1(g7573B));
AND2_X1 U_g3987B (.ZN(g3987B),.A2(FE_OFN359_g18B),.A1(g243B));
AND2_X1 U_g4765B (.ZN(g4765B),.A2(FE_OFN307_g4010B),.A1(g491B));
AND2_X1 U_g11555B (.ZN(g11555B),.A2(FE_OFN27_g11519B),.A1(FE_OFN238_g1781B));
AND2_X1 U_g9857B (.ZN(g9857B),.A2(g9569B),.A1(g9734B));
AND2_X1 U_g8728B (.ZN(g8728B),.A2(g7915B),.A1(g8226B));
AND2_X1 U_g8730B (.ZN(g8730B),.A2(g7917B),.A1(g8230B));
AND2_X1 U_g8185B (.ZN(g8185B),.A2(g8234B),.A1(g664B));
AND2_X1 U_g5194B (.ZN(g5194B),.A2(FE_OFN299_g4457B),.A1(g1610B));
AND2_X1 U_g8385B (.ZN(g8385B),.A2(g8234B),.A1(g5255B));
AND2_X1 U_g4610B (.ZN(g4610B),.A2(g2212B),.A1(g3804B));
AND2_X1 U_g7902B (.ZN(g7902B),.A2(g6449B),.A1(g7661B));
AND2_X1 U_g4073B (.ZN(g4073B),.A2(g3222B),.A1(g3200B));
AND2_X1 U_g8070B (.ZN(g8070B),.A2(FE_OFN198_g7697B),.A1(g682B));
AND2_X1 U_g5731B (.ZN(g5731B),.A2(FE_OFN315_g5117B),.A1(g1583B));
AND2_X1 U_g11238B (.ZN(g11238B),.A2(g11111B),.A1(g4553B));
AND2_X1 U_g4473B (.ZN(g4473B),.A2(FE_OFN302_g3913B),.A1(g1125B));
AND2_X1 U_g8470B (.ZN(g8470B),.A2(FE_OFN210_g7246B),.A1(g8308B));
AND2_X1 U_g5489B (.ZN(g5489B),.A2(FE_OFN358_g3521B),.A1(g557B));
AND2_X1 U_g3991B (.ZN(g3991B),.A2(g2774B),.A1(g1738B));
AND4_X1 U_I5887B (.ZN(I5887B),.A4(g2095B),.A3(g166B),.A2(g2083B),.A1(g2078B));
AND2_X1 U_g7823B (.ZN(g7823B),.A2(FE_OFN209_g6863B),.A1(g1923B));
AND2_X1 U_g4069B (.ZN(g4069B),.A2(g2777B),.A1(g1762B));
AND3_X4 U_g11519B (.ZN(g11519B),.A3(g11492B),.A2(g3015B),.A1(g1317B));
AND2_X1 U_g11176B (.ZN(g11176B),.A2(FE_OFN20_g10702B),.A1(g506B));
AND2_X1 U_g11092B (.ZN(g11092B),.A2(FE_OFN4_g10950B),.A1(g837B));
AND2_X1 U_g11154B (.ZN(g11154B),.A2(FE_OFN278_g10927B),.A1(g330B));
AND2_X1 U_g9608B (.ZN(g9608B),.A2(FE_OFN71_g9292B),.A1(g7B));
AND2_X1 U_g11637B (.ZN(g11637B),.A2(FE_OFN99_g4421B),.A1(g11596B));
AND2_X1 U_g2091B (.ZN(g2091B),.A2(g971B),.A1(g976B));
AND2_X1 U_g8406B (.ZN(g8406B),.A2(g8146B),.A1(g695B));
AND2_X1 U_g5254B (.ZN(g5254B),.A2(FE_OFN357_g3521B),.A1(g549B));
AND2_X1 U_g7260B (.ZN(g7260B),.A2(g2345B),.A1(g6752B));
AND2_X1 U_g5150B (.ZN(g5150B),.A2(g4678B),.A1(g1275B));
AND2_X1 U_g8766B (.ZN(g8766B),.A2(FE_OFN304_g5151B),.A1(g8612B));
AND2_X1 U_g9588B (.ZN(g9588B),.A2(FE_OFN53_g9173B),.A1(g1351B));
AND2_X1 U_g8801B (.ZN(g8801B),.A2(FE_OFN331_g8696B),.A1(g8742B));
AND2_X1 U_g7063B (.ZN(g7063B),.A2(g6586B),.A1(g5008B));
AND2_X1 U_g10303B (.ZN(g10303B),.A2(g9291B),.A1(g9995B));
AND2_X1 U_g5009B (.ZN(g5009B),.A2(FE_OFN154_g4640B),.A1(g1486B));
AND2_X1 U_g9665B (.ZN(g9665B),.A2(FE_OFN48_g9151B),.A1(g1314B));
AND2_X2 U_g8748B (.ZN(g8748B),.A2(g8488B),.A1(I9810B));
AND2_X1 U_g11215B (.ZN(g11215B),.A2(FE_OFN279_g11157B),.A1(g953B));
AND2_X1 U_g10750B (.ZN(g10750B),.A2(FE_OFN102_g3586B),.A1(g10597B));
AND3_X1 U_g5769B (.ZN(g5769B),.A3(g3818B),.A2(FE_OFN200_g4921B),.A1(g3092B));
AND2_X1 U_g6673B (.ZN(g6673B),.A2(I9326B),.A1(g90B));
AND2_X1 U_g5212B (.ZN(g5212B),.A2(g4678B),.A1(g1255B));
AND2_X1 U_g7720B (.ZN(g7720B),.A2(FE_OFN191_g6488B),.A1(g727B));
AND3_X1 U_g5918B (.ZN(g5918B),.A3(g4609B),.A2(FE_OFN184_I7048B),.A1(g109B));
AND2_X1 U_g8045B (.ZN(g8045B),.A2(g5128B),.A1(g7547B));
AND2_X1 U_g8173B (.ZN(g8173B),.A2(FE_OFN363_I5565B),.A1(g7971B));
AND2_X1 U_g11349B (.ZN(g11349B),.A2(g7914B),.A1(g11288B));
AND2_X1 U_g7843B (.ZN(g7843B),.A2(g5919B),.A1(g7599B));
AND2_X1 U_g9696B (.ZN(g9696B),.A2(FE_OFN59_g9432B),.A1(g281B));
AND2_X1 U_g6772B (.ZN(g6772B),.A2(g722B),.A1(g6228B));
AND2_X1 U_g6058B (.ZN(g6058B),.A2(g85B),.A1(g1035B));
AND2_X1 U_g6531B (.ZN(g6531B),.A2(FE_OFN283_I8869B),.A1(g79B));
AND2_X1 U_g6743B (.ZN(g6743B),.A2(FE_OFN219_g5557B),.A1(g4106B));
AND2_X1 U_g6890B (.ZN(g6890B),.A2(g6403B),.A1(g6752B));
AND2_X1 U_g7549B (.ZN(g7549B),.A2(FE_OFN137_g3829B),.A1(g7269B));
AND2_X1 U_g8169B (.ZN(g8169B),.A2(I11360B),.A1(g35B));
AND2_X1 U_g11304B (.ZN(g11304B),.A2(g11243B),.A1(g4585B));
AND2_X1 U_g9944B (.ZN(g9944B),.A2(FE_OFN68_g9392B),.A1(g9924B));
AND2_X4 U_g9240B (.ZN(g9240B),.A2(g8962B),.A1(FE_OFN277_g48B));
AND2_X1 U_g8059B (.ZN(g8059B),.A2(FE_OFN177_g5919B),.A1(g7592B));
AND2_X1 U_g8718B (.ZN(g8718B),.A2(g7903B),.A1(g8203B));
AND2_X1 U_g8767B (.ZN(g8767B),.A2(FE_OFN304_g5151B),.A1(g8616B));
AND2_X1 U_g9316B (.ZN(g9316B),.A2(g48B),.A1(g8877B));
AND2_X1 U_g7625B (.ZN(g7625B),.A2(FE_OFN191_g6488B),.A1(g673B));
AND2_X1 U_g8793B (.ZN(g8793B),.A2(FE_OFN331_g8696B),.A1(g8644B));
AND2_X1 U_g2940B (.ZN(g2940B),.A2(g1654B),.A1(g2424B));
AND2_X1 U_g4114B (.ZN(g4114B),.A2(g3301B),.A1(g1351B));
AND2_X1 U_g11636B (.ZN(g11636B),.A2(g7897B),.A1(g11624B));
AND2_X1 U_g10949B (.ZN(g10949B),.A2(g10809B),.A1(g2947B));
AND2_X1 U_g3563B (.ZN(g3563B),.A2(g2126B),.A1(g3275B));
AND2_X1 U_g10948B (.ZN(g10948B),.A2(g10809B),.A1(g2223B));
AND2_X1 U_g8246B (.ZN(g8246B),.A2(g7438B),.A1(g7846B));
AND2_X1 U_g5788B (.ZN(g5788B),.A2(g5222B),.A1(g1540B));
AND2_X1 U_g4008B (.ZN(g4008B),.A2(FE_OFN224_g2276B),.A1(FE_OFN236_g1776B));
AND2_X1 U_g9596B (.ZN(g9596B),.A2(g9010B),.A1(g928B));
AND2_X1 U_g5249B (.ZN(g5249B),.A2(FE_OFN288_g4263B),.A1(g1089B));
AND2_X1 U_g11585B (.ZN(g11585B),.A2(g11539B),.A1(g1321B));
AND2_X1 U_g3089B (.ZN(g3089B),.A2(g2050B),.A1(g2054B));
AND2_X1 U_g4972B (.ZN(g4972B),.A2(FE_OFN147_g4682B),.A1(g1436B));
AND2_X1 U_g11554B (.ZN(g11554B),.A2(FE_OFN27_g11519B),.A1(g1776B));
AND2_X1 U_g7586B (.ZN(g7586B),.A2(g5420B),.A1(g7096B));
AND2_X1 U_g10673B (.ZN(g10673B),.A2(FE_OFN79_g8700B),.A1(g10417B));
AND3_X1 U_g4806B (.ZN(g4806B),.A3(g2493B),.A2(g3992B),.A1(g3215B));
AND2_X1 U_g5485B (.ZN(g5485B),.A2(FE_OFN333_g4294B),.A1(g1914B));
AND2_X1 U_g9936B (.ZN(g9936B),.A2(FE_OFN60_g9624B),.A1(g9915B));
AND2_X1 U_g2910B (.ZN(g2910B),.A2(g1660B),.A1(g2424B));
AND2_X1 U_g9317B (.ZN(g9317B),.A2(g8875B),.A1(g6109B));
AND2_X1 U_g10933B (.ZN(g10933B),.A2(g3982B),.A1(g10853B));
AND2_X1 U_g8388B (.ZN(g8388B),.A2(g7246B),.A1(g8177B));
AND2_X1 U_g4465B (.ZN(g4465B),.A2(FE_OFN302_g3913B),.A1(g1117B));
AND2_X1 U_g7141B (.ZN(g7141B),.A2(g6716B),.A1(g5230B));
AND2_X1 U_g10508B (.ZN(g10508B),.A2(FE_OFN336_g1690B),.A1(g10013B));
AND2_X1 U_g4230B (.ZN(g4230B),.A2(FE_OFN132_g3015B),.A1(g1095B));
AND2_X1 U_g10634B (.ZN(g10634B),.A2(g3829B),.A1(g10382B));
AND2_X1 U_g9601B (.ZN(g9601B),.A2(g9192B),.A1(g922B));
AND2_X1 U_g6126B (.ZN(g6126B),.A2(FE_OFN322_g4449B),.A1(g3681B));
AND2_X1 U_g6326B (.ZN(g6326B),.A2(FE_OFN115_g4807B),.A1(g1250B));
AND2_X1 U_g7710B (.ZN(g7710B),.A2(FE_OFN191_g6488B),.A1(g700B));
AND2_X1 U_g8028B (.ZN(g8028B),.A2(g7438B),.A1(g7375B));
AND2_X1 U_g6760B (.ZN(g6760B),.A2(g6221B),.A1(g786B));
AND2_X1 U_g5640B (.ZN(g5640B),.A2(FE_OFN290_g4880B),.A1(g1059B));
AND2_X1 U_g5031B (.ZN(g5031B),.A2(FE_OFN153_g4640B),.A1(g1478B));
AND2_X1 U_g4550B (.ZN(g4550B),.A2(FE_OFN344_g3586B),.A1(g342B));
AND2_X1 U_g7879B (.ZN(g7879B),.A2(FE_OFN366_g3521B),.A1(g5286B));
AND2_X1 U_g7962B (.ZN(g7962B),.A2(g6403B),.A1(g7730B));
AND2_X1 U_g9597B (.ZN(g9597B),.A2(FE_OFN46_g9125B),.A1(g1170B));
AND2_X1 U_g10452B (.ZN(g10452B),.A2(FE_OFN234_g2024B),.A1(g10439B));
AND2_X1 U_g4891B (.ZN(g4891B),.A2(g4739B),.A1(g631B));
AND2_X1 U_g5005B (.ZN(g5005B),.A2(FE_OFN154_g4640B),.A1(g1490B));
AND2_X1 U_g6423B (.ZN(g6423B),.A2(FE_OFN217_g5013B),.A1(g4348B));
AND2_X1 U_g8108B (.ZN(g8108B),.A2(g7952B),.A1(g1891B));
AND3_X4 U_g4807B (.ZN(g4807B),.A3(I6360B),.A2(g1289B),.A1(g3015B));
AND2_X1 U_g5911B (.ZN(g5911B),.A2(g4977B),.A1(g3322B));
AND2_X1 U_g9937B (.ZN(g9937B),.A2(FE_OFN60_g9624B),.A1(g9916B));
AND2_X1 U_g9840B (.ZN(g9840B),.A2(g9747B),.A1(g9704B));
AND2_X1 U_g10780B (.ZN(g10780B),.A2(g4467B),.A1(g10723B));
AND2_X1 U_g8217B (.ZN(g8217B),.A2(g7883B),.A1(g1872B));
AND2_X1 U_g11013B (.ZN(g11013B),.A2(FE_OFN18_g10702B),.A1(g5209B));
AND2_X1 U_g9390B (.ZN(g9390B),.A2(FE_OFN48_g9151B),.A1(g1333B));
AND2_X1 U_g11214B (.ZN(g11214B),.A2(FE_OFN279_g11157B),.A1(g950B));
AND2_X1 U_g6327B (.ZN(g6327B),.A2(FE_OFN115_g4807B),.A1(g1255B));
AND2_X1 U_g4342B (.ZN(g4342B),.A2(FE_OFN351_g3913B),.A1(g1149B));
AND2_X1 U_g5796B (.ZN(g5796B),.A2(FE_OFN321_g5261B),.A1(g1564B));
AND2_X1 U_g5473B (.ZN(g5473B),.A2(FE_OFN367_g3521B),.A1(g546B));
AND2_X1 U_g6346B (.ZN(g6346B),.A2(g5878B),.A1(g5038B));
AND2_X1 U_g6633B (.ZN(g6633B),.A2(FE_OFN282_g6165B),.A1(g354B));
AND2_X1 U_g11005B (.ZN(g11005B),.A2(FE_OFN13_g10702B),.A1(g5119B));
AND2_X1 U_g8365B (.ZN(g8365B),.A2(g8146B),.A1(g668B));
AND2_X1 U_g8048B (.ZN(g8048B),.A2(g5919B),.A1(g7558B));
AND2_X1 U_g4481B (.ZN(g4481B),.A2(g3906B),.A1(g1713B));
AND2_X1 U_g4097B (.ZN(g4097B),.A2(g3060B),.A1(g2677B));
AND2_X1 U_g8055B (.ZN(g8055B),.A2(FE_OFN305_g5151B),.A1(g7588B));
AND2_X1 U_g4497B (.ZN(g4497B),.A2(FE_OFN344_g3586B),.A1(g351B));
AND2_X1 U_g9942B (.ZN(g9942B),.A2(FE_OFN67_g9367B),.A1(g9922B));
AND2_X1 U_g6696B (.ZN(g6696B),.A2(I9326B),.A1(g94B));
AND3_X1 U_g10731B (.ZN(g10731B),.A3(g10665B),.A2(g1850B),.A1(g5118B));
AND2_X1 U_g8827B (.ZN(g8827B),.A2(g8696B),.A1(g8552B));
AND2_X1 U_g5540B (.ZN(g5540B),.A2(g4292B),.A1(g1727B));
AND2_X1 U_g4960B (.ZN(g4960B),.A2(FE_OFN147_g4682B),.A1(g1403B));
AND2_X1 U_g8846B (.ZN(g8846B),.A2(FE_OFN328_g8709B),.A1(g8615B));
AND2_X1 U_g6508B (.ZN(g6508B),.A2(FE_OFN363_I5565B),.A1(g5983B));
AND2_X1 U_g6240B (.ZN(g6240B),.A2(g5361B),.A1(g182B));
AND2_X1 U_g7931B (.ZN(g7931B),.A2(g7446B),.A1(g52B));
AND2_X1 U_g5287B (.ZN(g5287B),.A2(g4782B),.A1(I6260B));
AND2_X1 U_g6472B (.ZN(g6472B),.A2(g1936B),.A1(g5853B));
AND2_X1 U_g11100B (.ZN(g11100B),.A2(FE_OFN4_g10950B),.A1(g853B));
AND2_X1 U_g11235B (.ZN(g11235B),.A2(g11107B),.A1(g4529B));
AND2_X1 U_g5199B (.ZN(g5199B),.A2(FE_OFN288_g4263B),.A1(g1068B));
AND2_X1 U_g6316B (.ZN(g6316B),.A2(FE_OFN117_g4807B),.A1(g1270B));
AND2_X1 U_g7515B (.ZN(g7515B),.A2(g70B),.A1(FE_OFN85_g2176B));
AND2_X1 U_g10583B (.ZN(g10583B),.A2(g10515B),.A1(g10518B));
AND2_X1 U_g5781B (.ZN(g5781B),.A2(g5222B),.A1(g1537B));
AND2_X1 U_g8018B (.ZN(g8018B),.A2(g7438B),.A1(g7742B));
AND2_X1 U_g4401B (.ZN(g4401B),.A2(g3772B),.A1(g1845B));
AND3_X1 U_g8994B (.ZN(g8994B),.A3(g8783B),.A2(FE_OFN92_g2216B),.A1(g8110B));
AND2_X1 U_g2950B (.ZN(g2950B),.A2(g1666B),.A1(g2424B));
AND2_X1 U_g5510B (.ZN(g5510B),.A2(g4289B),.A1(g1630B));
AND2_X1 U_g6347B (.ZN(g6347B),.A2(FE_OFN320_g5361B),.A1(g275B));
AND2_X1 U_g9357B (.ZN(g9357B),.A2(g9223B),.A1(g962B));
AND2_X1 U_g4828B (.ZN(g4828B),.A2(g695B),.A1(g4106B));
AND2_X1 U_g11407B (.ZN(g11407B),.A2(g4807B),.A1(g11249B));
AND2_X1 U_g4727B (.ZN(g4727B),.A2(FE_OFN300_g4002B),.A1(g386B));
AND2_X1 U_g10357B (.ZN(g10357B),.A2(FE_OFN269_g109B),.A1(I15500B));
AND2_X1 U_g10743B (.ZN(g10743B),.A2(FE_OFN364_g3015B),.A1(g10639B));
AND2_X1 U_g5259B (.ZN(g5259B),.A2(g4739B),.A1(g627B));
AND2_X1 U_g5694B (.ZN(g5694B),.A2(FE_OFN365_g5361B),.A1(g162B));
AND2_X1 U_g10769B (.ZN(g10769B),.A2(FE_OFN297_g3015B),.A1(g10652B));
AND2_X1 U_g11584B (.ZN(g11584B),.A2(g11539B),.A1(g1318B));
AND2_X1 U_g4932B (.ZN(g4932B),.A2(FE_OFN290_g4880B),.A1(g1065B));
AND2_X1 U_g10768B (.ZN(g10768B),.A2(FE_OFN293_g3015B),.A1(g10649B));
AND2_X1 U_g6820B (.ZN(g6820B),.A2(FE_OFN178_g5354B),.A1(g1362B));
AND2_X1 U_g4068B (.ZN(g4068B),.A2(FE_OFN224_g2276B),.A1(FE_OFN251_g1801B));
AND2_X1 U_g6317B (.ZN(g6317B),.A2(FE_OFN117_g4807B),.A1(g1304B));
AND2_X1 U_g5215B (.ZN(g5215B),.A2(g3275B),.A1(g4276B));
AND2_X1 U_g4576B (.ZN(g4576B),.A2(g4010B),.A1(g530B));
AND2_X1 U_g6775B (.ZN(g6775B),.A2(g6231B),.A1(g822B));
AND2_X4 U_g3829B (.ZN(g3829B),.A2(g1696B),.A1(g2028B));
AND2_X1 U_g10662B (.ZN(g10662B),.A2(g10396B),.A1(g8700B));
AND2_X1 U_g8101B (.ZN(g8101B),.A2(FE_OFN207_g6863B),.A1(g5484B));
AND2_X1 U_g5825B (.ZN(g5825B),.A2(g5318B),.A1(g3204B));
AND4_X1 U_I6310B (.ZN(I6310B),.A4(g2435B),.A3(g2421B),.A2(g2407B),.A1(g2396B));
AND2_X1 U_g7884B (.ZN(g7884B),.A2(FE_OFN334_g7045B),.A1(g7457B));
AND2_X1 U_g5008B (.ZN(g5008B),.A2(FE_OFN303_g4678B),.A1(g1292B));
AND2_X1 U_g3974B (.ZN(g3974B),.A2(FE_OFN260_g18B),.A1(g231B));
AND2_X1 U_g9949B (.ZN(g9949B),.A2(FE_OFN68_g9392B),.A1(g9929B));
AND2_X1 U_g2531B (.ZN(g2531B),.A2(g668B),.A1(g658B));
AND2_X2 U_g9292B (.ZN(g9292B),.A2(g48B),.A1(g8878B));
AND2_X1 U_g10778B (.ZN(g10778B),.A2(g10679B),.A1(g1027B));
AND2_X1 U_g8041B (.ZN(g8041B),.A2(g5128B),.A1(g7524B));
AND2_X1 U_g6079B (.ZN(g6079B),.A2(FE_OFN273_g85B),.A1(g1053B));
AND2_X1 U_g7235B (.ZN(g7235B),.A2(g6447B),.A1(g6663B));
AND2_X1 U_g9603B (.ZN(g9603B),.A2(FE_OFN46_g9125B),.A1(g1173B));
AND2_X1 U_g6840B (.ZN(g6840B),.A2(FE_OFN180_g5354B),.A1(g248B));
AND2_X1 U_g9850B (.ZN(g9850B),.A2(g9579B),.A1(g9726B));
AND2_X1 U_g7988B (.ZN(g7988B),.A2(g7379B),.A1(g1878B));
AND2_X1 U_g5228B (.ZN(g5228B),.A2(FE_OFN288_g4263B),.A1(g1086B));
AND2_X1 U_g7134B (.ZN(g7134B),.A2(g6354B),.A1(g5587B));
AND2_X1 U_g5934B (.ZN(g5934B),.A2(g1965B),.A1(g5215B));
AND2_X1 U_g5230B (.ZN(g5230B),.A2(g4678B),.A1(g1265B));
AND2_X1 U_g8168B (.ZN(g8168B),.A2(FE_OFN89_I11360B),.A1(g34B));
AND2_X1 U_g9583B (.ZN(g9583B),.A2(g8995B),.A1(g886B));
AND2_X1 U_g10672B (.ZN(g10672B),.A2(g9473B),.A1(g10414B));
AND2_X1 U_g3287B (.ZN(g3287B),.A2(g5188B),.A1(g802B));
AND2_X1 U_g8772B (.ZN(g8772B),.A2(FE_OFN304_g5151B),.A1(g8627B));
AND2_X1 U_g4893B (.ZN(g4893B),.A2(g4739B),.A1(g635B));
AND2_X1 U_g10331B (.ZN(g10331B),.A2(FE_OFN269_g109B),.A1(I15510B));
AND2_X1 U_g8505B (.ZN(g8505B),.A2(FE_OFN359_g18B),.A1(g8309B));
AND2_X1 U_g10449B (.ZN(g10449B),.A2(FE_OFN235_g2024B),.A1(g10433B));
AND2_X1 U_g11273B (.ZN(g11273B),.A2(g11199B),.A1(g4765B));
AND2_X1 U_g8734B (.ZN(g8734B),.A2(g7923B),.A1(g8187B));
AND2_X1 U_g5913B (.ZN(g5913B),.A2(g85B),.A1(g1041B));
AND2_X1 U_g10448B (.ZN(g10448B),.A2(FE_OFN235_g2024B),.A1(g10421B));
AND2_X1 U_g6163B (.ZN(g6163B),.A2(g5354B),.A1(g4572B));
AND2_X1 U_g6363B (.ZN(g6363B),.A2(FE_OFN320_g5361B),.A1(g284B));
AND2_X1 U_g7202B (.ZN(g7202B),.A2(FE_OFN322_g4449B),.A1(g5226B));
AND2_X1 U_g11463B (.ZN(g11463B),.A2(FE_OFN99_g4421B),.A1(g11229B));
AND2_X1 U_g8074B (.ZN(g8074B),.A2(FE_OFN198_g7697B),.A1(g718B));
AND2_X1 U_g4325B (.ZN(g4325B),.A2(FE_OFN351_g3913B),.A1(g1166B));
AND2_X1 U_g8474B (.ZN(g8474B),.A2(g5521B),.A1(g8383B));
AND2_X1 U_g11234B (.ZN(g11234B),.A2(g11107B),.A1(g4518B));
AND2_X1 U_g5266B (.ZN(g5266B),.A2(FE_OFN335_g4737B),.A1(g718B));
AND2_X1 U_g4483B (.ZN(g4483B),.A2(FE_OFN103_g3586B),.A1(g336B));
AND2_X1 U_g5248B (.ZN(g5248B),.A2(FE_OFN335_g4737B),.A1(g673B));
AND2_X1 U_g11514B (.ZN(g11514B),.A2(FE_OFN176_g5151B),.A1(g11491B));
AND2_X1 U_g5255B (.ZN(g5255B),.A2(FE_OFN335_g4737B),.A1(g682B));
AND2_X1 U_g4106B (.ZN(g4106B),.A2(g686B),.A1(g3284B));
AND2_X1 U_g2760B (.ZN(g2760B),.A2(g2091B),.A1(g981B));
AND2_X1 U_g5097B (.ZN(g5097B),.A2(g4608B),.A1(g1786B));
AND2_X1 U_g5726B (.ZN(g5726B),.A2(FE_OFN315_g5117B),.A1(g1601B));
AND2_X1 U_g5497B (.ZN(g5497B),.A2(FE_OFN357_g3521B),.A1(g560B));
AND2_X4 U_g5354B (.ZN(g5354B),.A2(I7048B),.A1(FE_OFN352_g109B));
AND2_X1 U_g7933B (.ZN(g7933B),.A2(g7450B),.A1(g55B));
AND2_X1 U_g9617B (.ZN(g9617B),.A2(g9274B),.A1(g9B));
AND2_X1 U_g9906B (.ZN(g9906B),.A2(g9680B),.A1(g9873B));
AND2_X1 U_g11012B (.ZN(g11012B),.A2(FE_OFN18_g10702B),.A1(g5196B));
AND2_X1 U_g7050B (.ZN(g7050B),.A2(g6702B),.A1(g5001B));
AND2_X1 U_g10971B (.ZN(g10971B),.A2(g2045B),.A1(g10849B));
AND2_X1 U_g4904B (.ZN(g4904B),.A2(g4243B),.A1(g1850B));
AND2_X1 U_g10369B (.ZN(g10369B),.A2(FE_OFN235_g2024B),.A1(g10361B));
AND2_X1 U_g8400B (.ZN(g8400B),.A2(g8234B),.A1(g5271B));
AND2_X1 U_g4345B (.ZN(g4345B),.A2(FE_OFN289_g4679B),.A1(g1169B));
AND2_X1 U_g2161B (.ZN(g2161B),.A2(I5085B),.A1(I5084B));
AND2_X1 U_g5001B (.ZN(g5001B),.A2(FE_OFN303_g4678B),.A1(g1300B));
AND2_X1 U_g9945B (.ZN(g9945B),.A2(FE_OFN68_g9392B),.A1(g9925B));
AND2_X1 U_g7271B (.ZN(g7271B),.A2(g6354B),.A1(g5028B));
AND2_X1 U_g9709B (.ZN(g9709B),.A2(FE_OFN70_g9490B),.A1(g1524B));
AND2_X1 U_g4223B (.ZN(g4223B),.A2(FE_OFN347_g3914B),.A1(g1003B));
AND2_X1 U_g10716B (.ZN(g10716B),.A2(g10396B),.A1(g10497B));
AND2_X1 U_g11291B (.ZN(g11291B),.A2(g4379B),.A1(g11247B));
AND2_X1 U_g6661B (.ZN(g6661B),.A2(FE_OFN97_I8869B),.A1(g73B));
AND2_X1 U_g11173B (.ZN(g11173B),.A2(FE_OFN21_g10702B),.A1(g491B));
AND2_X1 U_g6075B (.ZN(g6075B),.A2(g5613B),.A1(g549B));
AND2_X1 U_g8023B (.ZN(g8023B),.A2(g7438B),.A1(g7367B));
AND2_X1 U_g9907B (.ZN(g9907B),.A2(g9680B),.A1(g9888B));
AND2_X1 U_g10582B (.ZN(g10582B),.A2(g9473B),.A1(g10339B));
AND2_X1 U_g5746B (.ZN(g5746B),.A2(FE_OFN353_g5117B),.A1(g1589B));
AND2_X1 U_g5221B (.ZN(g5221B),.A2(g4678B),.A1(g1260B));
AND2_X1 U_g9959B (.ZN(g9959B),.A2(FE_OFN280_g9536B),.A1(g9950B));
AND2_X1 U_g7674B (.ZN(g7674B),.A2(g3880B),.A1(g5857B));
AND2_X1 U_g9690B (.ZN(g9690B),.A2(g9432B),.A1(g266B));
AND2_X1 U_g6627B (.ZN(g6627B),.A2(FE_OFN283_I8869B),.A1(g58B));
AND2_X1 U_g5703B (.ZN(g5703B),.A2(FE_OFN365_g5361B),.A1(g174B));
AND2_X1 U_g4522B (.ZN(g4522B),.A2(FE_OFN344_g3586B),.A1(g360B));
AND2_X1 U_g4115B (.ZN(g4115B),.A2(g3060B),.A1(FE_OFN236_g1776B));
AND2_X1 U_g7541B (.ZN(g7541B),.A2(I6360B),.A1(g7075B));
AND2_X1 U_g10627B (.ZN(g10627B),.A2(FE_OFN227_g3880B),.A1(g10452B));
AND2_X1 U_g4047B (.ZN(g4047B),.A2(FE_OFN225_g2276B),.A1(FE_OFN238_g1781B));
AND2_X1 U_g6526B (.ZN(g6526B),.A2(FE_OFN283_I8869B),.A1(g76B));
AND2_X1 U_g2944B (.ZN(g2944B),.A2(g1669B),.A1(g2424B));
AND2_X1 U_g6646B (.ZN(g6646B),.A2(g6165B),.A1(g360B));
AND2_X1 U_g7132B (.ZN(g7132B),.A2(g6702B),.A1(g5182B));
AND2_X1 U_g11029B (.ZN(g11029B),.A2(FE_OFN17_g10702B),.A1(g401B));
AND2_X1 U_g8051B (.ZN(g8051B),.A2(FE_OFN305_g5151B),.A1(g7572B));
AND2_X1 U_g8127B (.ZN(g8127B),.A2(g7949B),.A1(g1927B));
AND2_X1 U_g7209B (.ZN(g7209B),.A2(g6432B),.A1(g3804B));
AND2_X1 U_g11028B (.ZN(g11028B),.A2(FE_OFN17_g10702B),.A1(g396B));
AND2_X1 U_g6439B (.ZN(g6439B),.A2(g5919B),.A1(g3631B));
AND2_X1 U_g10742B (.ZN(g10742B),.A2(g3586B),.A1(g10655B));
AND2_X1 U_g9110B (.ZN(g9110B),.A2(FE_OFN359_g18B),.A1(g8880B));
AND2_X1 U_g10681B (.ZN(g10681B),.A2(g3586B),.A1(g10567B));
AND2_X1 U_g4537B (.ZN(g4537B),.A2(g4002B),.A1(g444B));
AND2_X1 U_g9663B (.ZN(g9663B),.A2(FE_OFN39_g9223B),.A1(g959B));
AND2_X1 U_g5349B (.ZN(g5349B),.A2(g4617B),.A1(g2126B));
AND2_X1 U_g8732B (.ZN(g8732B),.A2(g7919B),.A1(g8200B));
AND2_X1 U_g3807B (.ZN(g3807B),.A2(g3062B),.A1(g3003B));
AND2_X1 U_g5848B (.ZN(g5848B),.A2(g5519B),.A1(g3860B));
AND2_X1 U_g8508B (.ZN(g8508B),.A2(FE_OFN330_g7638B),.A1(g8411B));
AND2_X1 U_g8072B (.ZN(g8072B),.A2(FE_OFN199_g7697B),.A1(g700B));
AND2_X1 U_g5699B (.ZN(g5699B),.A2(g5117B),.A1(g1592B));
AND2_X1 U_g11240B (.ZN(g11240B),.A2(g11111B),.A1(g4560B));
AND2_X1 U_g5398B (.ZN(g5398B),.A2(g2224B),.A1(g4610B));
AND2_X1 U_g6616B (.ZN(g6616B),.A2(FE_OFN363_I5565B),.A1(g6105B));
AND2_X1 U_g10690B (.ZN(g10690B),.A2(FE_OFN136_g3863B),.A1(g10387B));
AND2_X1 U_g8043B (.ZN(g8043B),.A2(FE_OFN305_g5151B),.A1(g7582B));
AND2_X1 U_g9590B (.ZN(g9590B),.A2(g8995B),.A1(g895B));
AND2_X1 U_g4128B (.ZN(g4128B),.A2(g627B),.A1(g1976B));
AND2_X1 U_g6404B (.ZN(g6404B),.A2(FE_OFN217_g5013B),.A1(g2132B));
AND2_X1 U_g6647B (.ZN(g6647B),.A2(g5808B),.A1(g87B));
AND2_X1 U_g10504B (.ZN(g10504B),.A2(FE_OFN336_g1690B),.A1(g10001B));
AND2_X1 U_g9657B (.ZN(g9657B),.A2(g9205B),.A1(g919B));
AND2_X1 U_g4542B (.ZN(g4542B),.A2(FE_OFN344_g3586B),.A1(g366B));
AND2_X1 U_g4330B (.ZN(g4330B),.A2(FE_OFN351_g3913B),.A1(g1163B));
AND2_X1 U_g3497B (.ZN(g3497B),.A2(g1900B),.A1(g2804B));
AND2_X1 U_g5524B (.ZN(g5524B),.A2(g3906B),.A1(g1678B));
AND2_X1 U_g8147B (.ZN(g8147B),.A2(g7907B),.A1(g928B));
AND2_X1 U_g4554B (.ZN(g4554B),.A2(g4010B),.A1(g542B));
AND2_X1 U_g9899B (.ZN(g9899B),.A2(g9367B),.A1(g9713B));
AND2_X1 U_g5258B (.ZN(g5258B),.A2(FE_OFN335_g4737B),.A1(g700B));
AND2_X1 U_g7736B (.ZN(g7736B),.A2(FE_OFN226_g3880B),.A1(g5814B));
AND2_X1 U_g6224B (.ZN(g6224B),.A2(FE_OFN306_g5128B),.A1(g1520B));
AND2_X1 U_g10626B (.ZN(g10626B),.A2(FE_OFN369_g4525B),.A1(g10453B));
AND2_X1 U_g6320B (.ZN(g6320B),.A2(FE_OFN118_g4807B),.A1(g1292B));
AND2_X1 U_g7623B (.ZN(g7623B),.A2(FE_OFN191_g6488B),.A1(g664B));
AND2_X1 U_g10299B (.ZN(g10299B),.A2(g10013B),.A1(FE_OFN76_g8700B));
AND2_X1 U_g7889B (.ZN(g7889B),.A2(g3814B),.A1(g5304B));
AND2_X1 U_g10298B (.ZN(g10298B),.A2(g10007B),.A1(g8700B));
AND2_X1 U_g8413B (.ZN(g8413B),.A2(g8146B),.A1(g722B));
AND2_X1 U_g3979B (.ZN(g3979B),.A2(FE_OFN260_g18B),.A1(g237B));
AND2_X1 U_g4902B (.ZN(g4902B),.A2(g4243B),.A1(g1848B));
AND2_X1 U_g5211B (.ZN(g5211B),.A2(FE_OFN288_g4263B),.A1(g1080B));
AND2_X1 U_g4512B (.ZN(g4512B),.A2(FE_OFN344_g3586B),.A1(g357B));
AND2_X1 U_g7722B (.ZN(g7722B),.A2(g6449B),.A1(g7127B));
AND2_X1 U_g9844B (.ZN(g9844B),.A2(g9522B),.A1(g9714B));
AND2_X1 U_g4490B (.ZN(g4490B),.A2(FE_OFN302_g3913B),.A1(g1141B));
AND2_X1 U_g6516B (.ZN(g6516B),.A2(FE_OFN363_I5565B),.A1(g5993B));
AND2_X1 U_g5026B (.ZN(g5026B),.A2(FE_OFN153_g4640B),.A1(g1453B));
AND2_X1 U_g8820B (.ZN(g8820B),.A2(g4737B),.A1(g8705B));
AND2_X1 U_g10737B (.ZN(g10737B),.A2(FE_OFN133_g3015B),.A1(g10597B));
AND3_X1 U_g8936B (.ZN(g8936B),.A3(g8849B),.A2(FE_OFN93_g2216B),.A1(g8115B));
AND2_X1 U_g10232B (.ZN(g10232B),.A2(g9974B),.A1(FE_OFN76_g8700B));
AND2_X1 U_g6771B (.ZN(g6771B),.A2(FE_OFN320_g5361B),.A1(g263B));
AND2_X1 U_g5170B (.ZN(g5170B),.A2(g4457B),.A1(g1811B));
AND2_X1 U_g8117B (.ZN(g8117B),.A2(FE_OFN207_g6863B),.A1(g5514B));
AND2_X1 U_g4529B (.ZN(g4529B),.A2(g4002B),.A1(g448B));
AND2_X1 U_g4348B (.ZN(g4348B),.A2(g1909B),.A1(g3497B));
AND2_X1 U_g9966B (.ZN(g9966B),.A2(FE_OFN280_g9536B),.A1(g9956B));
AND2_X1 U_g5280B (.ZN(g5280B),.A2(g2118B),.A1(g3967B));
AND2_X1 U_g7139B (.ZN(g7139B),.A2(g6716B),.A1(g5212B));
AND2_X1 U_g11099B (.ZN(g11099B),.A2(g10883B),.A1(g382B));
AND2_X1 U_g6892B (.ZN(g6892B),.A2(g5013B),.A1(g6472B));
AND2_X1 U_g9705B (.ZN(g9705B),.A2(g9474B),.A1(g1580B));
AND2_X1 U_g10512B (.ZN(g10512B),.A2(FE_OFN336_g1690B),.A1(g10025B));
AND2_X1 U_g11098B (.ZN(g11098B),.A2(FE_OFN4_g10950B),.A1(g849B));
AND2_X1 U_g8775B (.ZN(g8775B),.A2(FE_OFN304_g5151B),.A1(g8628B));
AND2_X1 U_g5083B (.ZN(g5083B),.A2(g4782B),.A1(g2510B));
AND2_X1 U_g5544B (.ZN(g5544B),.A2(FE_OFN291_g4880B),.A1(g1687B));
AND2_X1 U_g11272B (.ZN(g11272B),.A2(g11199B),.A1(g4760B));
AND2_X1 U_g5483B (.ZN(g5483B),.A2(g3906B),.A1(g1621B));
AND2_X1 U_g9948B (.ZN(g9948B),.A2(FE_OFN68_g9392B),.A1(g9928B));
AND2_X1 U_g4063B (.ZN(g4063B),.A2(FE_OFN224_g2276B),.A1(FE_OFN239_g1796B));
AND2_X1 U_g11462B (.ZN(g11462B),.A2(FE_OFN99_g4421B),.A1(g11227B));
AND2_X1 U_g6738B (.ZN(g6738B),.A2(FE_OFN219_g5557B),.A1(g2531B));
AND2_X1 U_g8060B (.ZN(g8060B),.A2(FE_OFN177_g5919B),.A1(g7593B));
AND2_X1 U_g6244B (.ZN(g6244B),.A2(FE_OFN306_g5128B),.A1(g1411B));
AND2_X1 U_g11032B (.ZN(g11032B),.A2(FE_OFN14_g10702B),.A1(g416B));
AND2_X1 U_g10445B (.ZN(g10445B),.A2(g1690B),.A1(g9974B));
AND2_X1 U_g9150B (.ZN(g9150B),.A2(FE_OFN325_g18B),.A1(g8882B));
AND2_X1 U_g10316B (.ZN(g10316B),.A2(g9097B),.A1(g10025B));
AND2_X1 U_g5756B (.ZN(g5756B),.A2(g5261B),.A1(g1531B));
AND2_X1 U_g4720B (.ZN(g4720B),.A2(g4673B),.A1(g1023B));
AND2_X1 U_g9409B (.ZN(g9409B),.A2(g9052B),.A1(g1721B));
AND2_X4 U_g8995B (.ZN(g8995B),.A2(g8929B),.A1(FE_OFN277_g48B));
AND2_X1 U_g6876B (.ZN(g6876B),.A2(g6557B),.A1(g4070B));
AND2_X1 U_g4989B (.ZN(g4989B),.A2(FE_OFN146_g4682B),.A1(g1424B));
AND2_X1 U_g9836B (.ZN(g9836B),.A2(FE_OFN34_g9785B),.A1(g9737B));
AND3_X1 U_g6656B (.ZN(g6656B),.A3(FE_OFN184_I7048B),.A2(g6061B),.A1(g109B));
AND2_X1 U_g5514B (.ZN(g5514B),.A2(FE_OFN333_g4294B),.A1(g1941B));
AND2_X1 U_g8390B (.ZN(g8390B),.A2(g6465B),.A1(g8268B));
AND2_X1 U_g5003B (.ZN(g5003B),.A2(FE_OFN154_g4640B),.A1(g1466B));
AND2_X1 U_g9967B (.ZN(g9967B),.A2(FE_OFN280_g9536B),.A1(g9957B));
AND2_X1 U_g5145B (.ZN(g5145B),.A2(g4673B),.A1(g1639B));
AND2_X1 U_g4971B (.ZN(g4971B),.A2(FE_OFN146_g4682B),.A1(g1419B));
AND2_X1 U_g10753B (.ZN(g10753B),.A2(FE_OFN133_g3015B),.A1(g10649B));
AND2_X1 U_g5695B (.ZN(g5695B),.A2(FE_OFN356_g5361B),.A1(g166B));
AND2_X1 U_g7613B (.ZN(g7613B),.A2(g5013B),.A1(g6940B));
AND2_X1 U_g10736B (.ZN(g10736B),.A2(FE_OFN293_g3015B),.A1(g10658B));
AND2_X1 U_g11220B (.ZN(g11220B),.A2(FE_OFN279_g11157B),.A1(g962B));
AND2_X1 U_g7444B (.ZN(g7444B),.A2(g5557B),.A1(g7277B));
AND2_X1 U_g5536B (.ZN(g5536B),.A2(FE_OFN310_g4336B),.A1(g2970B));
AND2_X1 U_g6663B (.ZN(g6663B),.A2(g2237B),.A1(g6064B));
AND2_X1 U_g4670B (.ZN(g4670B),.A2(g2355B),.A1(g192B));
AND2_X1 U_g6824B (.ZN(g6824B),.A2(FE_OFN178_g5354B),.A1(g1371B));
AND2_X1 U_g4253B (.ZN(g4253B),.A2(FE_OFN132_g3015B),.A1(g1074B));
AND2_X1 U_g8250B (.ZN(g8250B),.A2(g7907B),.A1(g932B));
AND2_X1 U_g8163B (.ZN(g8163B),.A2(g3737B),.A1(g7960B));
AND2_X1 U_g10764B (.ZN(g10764B),.A2(FE_OFN345_g3015B),.A1(g10643B));
AND2_X1 U_g5757B (.ZN(g5757B),.A2(g5222B),.A1(g1552B));
AND2_X1 U_g8032B (.ZN(g8032B),.A2(g7438B),.A1(g7385B));
AND2_X1 U_g11591B (.ZN(g11591B),.A2(g11561B),.A1(g2988B));
AND2_X1 U_g8053B (.ZN(g8053B),.A2(FE_OFN177_g5919B),.A1(g7583B));
AND2_X1 U_g11147B (.ZN(g11147B),.A2(FE_OFN278_g10927B),.A1(g321B));
AND2_X1 U_g5522B (.ZN(g5522B),.A2(g4289B),.A1(g1633B));
AND2_X1 U_g5115B (.ZN(g5115B),.A2(g4572B),.A1(g1394B));
AND2_X1 U_g9837B (.ZN(g9837B),.A2(g9751B),.A1(g9697B));
AND2_X1 U_g9620B (.ZN(g9620B),.A2(FE_OFN40_g9240B),.A1(g976B));
AND2_X1 U_g11151B (.ZN(g11151B),.A2(FE_OFN278_g10927B),.A1(g327B));
AND2_X1 U_g11172B (.ZN(g11172B),.A2(FE_OFN21_g10702B),.A1(g486B));
AND2_X1 U_g7885B (.ZN(g7885B),.A2(g3814B),.A1(g5300B));
AND2_X1 U_g6064B (.ZN(g6064B),.A2(g2230B),.A1(g5398B));
AND3_X1 U_g8929B (.ZN(g8929B),.A3(g8828B),.A2(FE_OFN95_g2216B),.A1(g8095B));
AND2_X1 U_g5595B (.ZN(g5595B),.A2(FE_OFN367_g3521B),.A1(g1621B));
AND2_X1 U_g5537B (.ZN(g5537B),.A2(g4449B),.A1(g2260B));
AND2_X1 U_g9842B (.ZN(g9842B),.A2(g9516B),.A1(g9708B));
AND2_X1 U_g4141B (.ZN(g4141B),.A2(g3060B),.A1(FE_OFN252_g1791B));
AND2_X1 U_g4341B (.ZN(g4341B),.A2(FE_OFN103_g3586B),.A1(g339B));
AND2_X4 U_g9192B (.ZN(g9192B),.A2(g8955B),.A1(FE_OFN277_g48B));
AND2_X1 U_g7679B (.ZN(g7679B),.A2(g6863B),.A1(g1950B));
AND2_X1 U_g7378B (.ZN(g7378B),.A2(FE_OFN226_g3880B),.A1(g5847B));
AND2_X1 U_g5612B (.ZN(g5612B),.A2(FE_OFN357_g3521B),.A1(g1627B));
AND2_X1 U_g7135B (.ZN(g7135B),.A2(g6355B),.A1(g869B));
AND2_X1 U_g10970B (.ZN(g10970B),.A2(g3390B),.A1(g10852B));
AND2_X1 U_g11025B (.ZN(g11025B),.A2(FE_OFN9_g10702B),.A1(g426B));
AND2_X1 U_g9854B (.ZN(g9854B),.A2(g9563B),.A1(g9730B));
AND2_X1 U_g7182B (.ZN(g7182B),.A2(FE_OFN213_g6003B),.A1(g1878B));
AND2_X1 U_g9941B (.ZN(g9941B),.A2(FE_OFN67_g9367B),.A1(g9921B));
AND2_X1 U_g6194B (.ZN(g6194B),.A2(FE_OFN289_g4679B),.A1(g554B));
AND2_X2 U_g5128B (.ZN(g5128B),.A2(FE_OFN352_g109B),.A1(I7048B));
AND2_X1 U_g4962B (.ZN(g4962B),.A2(g4467B),.A1(g1651B));
AND2_X1 U_g4358B (.ZN(g4358B),.A2(g3906B),.A1(g1209B));
AND2_X1 U_g8683B (.ZN(g8683B),.A2(g8549B),.A1(g4803B));
AND2_X1 U_g4506B (.ZN(g4506B),.A2(FE_OFN351_g3913B),.A1(g1113B));
AND2_X1 U_g6471B (.ZN(g6471B),.A2(g5878B),.A1(g5224B));
AND2_X1 U_g8778B (.ZN(g8778B),.A2(g1975B),.A1(g8688B));
AND2_X1 U_g11281B (.ZN(g11281B),.A2(g11203B),.A1(g4788B));
AND2_X1 U_g11146B (.ZN(g11146B),.A2(FE_OFN278_g10927B),.A1(g318B));
AND2_X1 U_g3904B (.ZN(g3904B),.A2(g627B),.A1(g2948B));
AND2_X1 U_g8075B (.ZN(g8075B),.A2(g7697B),.A1(g727B));
AND2_X1 U_g9829B (.ZN(g9829B),.A2(FE_OFN34_g9785B),.A1(g9723B));
AND3_X1 U_g8949B (.ZN(g8949B),.A3(g8828B),.A2(FE_OFN92_g2216B),.A1(g8255B));
AND2_X1 U_g7632B (.ZN(g7632B),.A2(g5420B),.A1(g7184B));
AND2_X1 U_g11290B (.ZN(g11290B),.A2(g4379B),.A1(g11246B));
AND2_X1 U_g6350B (.ZN(g6350B),.A2(FE_OFN346_g4381B),.A1(g5837B));
AND2_X1 U_g10599B (.ZN(g10599B),.A2(g4365B),.A1(g10448B));
AND2_X1 U_g5902B (.ZN(g5902B),.A2(g4977B),.A1(g2555B));
AND4_X1 U_I6337B (.ZN(I6337B),.A4(g2396B),.A3(g2407B),.A2(g2421B),.A1(g201B));
AND2_X2 U_g2276B (.ZN(g2276B),.A2(g1610B),.A1(g1765B));
AND2_X1 U_g6438B (.ZN(g6438B),.A2(g5013B),.A1(g5853B));
AND2_X1 U_g5512B (.ZN(g5512B),.A2(g4281B),.A1(g1660B));
AND2_X1 U_g5090B (.ZN(g5090B),.A2(FE_OFN299_g4457B),.A1(g1781B));
AND2_X1 U_g7719B (.ZN(g7719B),.A2(FE_OFN191_g6488B),.A1(g718B));
AND2_X1 U_g2561B (.ZN(g2561B),.A2(g741B),.A1(g742B));
AND2_X1 U_g3695B (.ZN(g3695B),.A2(FE_OFN292_g3015B),.A1(g1712B));
AND2_X1 U_g8603B (.ZN(g8603B),.A2(g8548B),.A1(g3983B));
AND2_X1 U_g8039B (.ZN(g8039B),.A2(FE_OFN305_g5151B),.A1(g7587B));
AND2_X1 U_g9610B (.ZN(g9610B),.A2(g9192B),.A1(g925B));
AND2_X1 U_g3536B (.ZN(g3536B),.A2(g3103B),.A1(g1289B));
AND2_X1 U_g5529B (.ZN(g5529B),.A2(FE_OFN310_g4336B),.A1(g2257B));
AND2_X1 U_g5148B (.ZN(g5148B),.A2(g4671B),.A1(g1107B));
AND2_X1 U_g9124B (.ZN(g9124B),.A2(FE_OFN325_g18B),.A1(g8881B));
AND2_X1 U_g9324B (.ZN(g9324B),.A2(FE_OFN275_g48B),.A1(g8879B));
AND2_X1 U_g4559B (.ZN(g4559B),.A2(FE_OFN137_g3829B),.A1(g2034B));
AND2_X1 U_g10561B (.ZN(g10561B),.A2(FE_OFN370_g4525B),.A1(g10549B));
AND2_X1 U_g5698B (.ZN(g5698B),.A2(FE_OFN315_g5117B),.A1(g1571B));
AND2_X1 U_g11226B (.ZN(g11226B),.A2(g11060B),.A1(g461B));
AND2_X1 U_g10295B (.ZN(g10295B),.A2(g9995B),.A1(FE_OFN79_g8700B));
AND2_X1 U_g5260B (.ZN(g5260B),.A2(FE_OFN288_g4263B),.A1(g1092B));
AND2_X1 U_g10680B (.ZN(g10680B),.A2(FE_OFN102_g3586B),.A1(g10564B));
AND2_X1 U_g6822B (.ZN(g6822B),.A2(FE_OFN178_g5354B),.A1(g231B));
AND2_X1 U_g4905B (.ZN(g4905B),.A2(g4243B),.A1(g1853B));
AND2_X1 U_g11551B (.ZN(g11551B),.A2(FE_OFN119_g3015B),.A1(g11538B));
AND2_X1 U_g3047B (.ZN(g3047B),.A2(g2306B),.A1(g1227B));
AND2_X1 U_g9849B (.ZN(g9849B),.A2(g9764B),.A1(g293B));
AND2_X1 U_g5279B (.ZN(g5279B),.A2(FE_OFN299_g4457B),.A1(g1766B));
AND2_X1 U_g8404B (.ZN(g8404B),.A2(g8146B),.A1(g686B));
AND2_X1 U_g5720B (.ZN(g5720B),.A2(FE_OFN168_g5361B),.A1(g170B));
AND2_X1 U_g5318B (.ZN(g5318B),.A2(g1857B),.A1(FE_OFN223_g4401B));
AND2_X1 U_g11376B (.ZN(g11376B),.A2(g4285B),.A1(g11318B));
AND2_X1 U_g11297B (.ZN(g11297B),.A2(g11243B),.A1(g4565B));
AND2_X1 U_g9898B (.ZN(g9898B),.A2(g9367B),.A1(g9710B));
OR2_X1 U_g6895B (.ZN(g6895B),.A2(g4875B),.A1(g6776B));
OR2_X1 U_g7189B (.ZN(g7189B),.A2(I9717B),.A1(g6632B));
OR2_X1 U_g9510B (.ZN(g9510B),.A2(g9111B),.A1(FE_OFN44_g9125B));
OR2_X1 U_g7297B (.ZN(g7297B),.A2(g6323B),.A1(g7132B));
OR2_X1 U_g9088B (.ZN(g9088B),.A2(g8233B),.A1(g8927B));
OR2_X1 U_g9923B (.ZN(g9923B),.A2(g9707B),.A1(g9865B));
OR2_X1 U_g6485B (.ZN(g6485B),.A2(g5067B),.A1(g5848B));
OR2_X1 U_g8771B (.ZN(g8771B),.A2(g8652B),.A1(g5483B));
OR2_X1 U_g5813B (.ZN(g5813B),.A2(g4869B),.A1(g5617B));
OR2_X1 U_g7963B (.ZN(g7963B),.A2(g7182B),.A1(FE_OFN334_g7045B));
OR2_X1 U_g10643B (.ZN(g10643B),.A2(g7736B),.A1(g10624B));
OR3_X1 U_g9886B (.ZN(g9886B),.A3(g9759B),.A2(g9592B),.A1(g9607B));
OR3_X1 U_g9951B (.ZN(g9951B),.A3(g9803B),.A2(g9899B),.A1(g9902B));
OR2_X1 U_g11625B (.ZN(g11625B),.A2(g11597B),.A1(g6535B));
OR2_X1 U_g8945B (.ZN(g8945B),.A2(FE_OFN332_g8748B),.A1(g8801B));
OR2_X1 U_g10489B (.ZN(g10489B),.A2(g10367B),.A1(g4456B));
OR2_X1 U_g10559B (.ZN(g10559B),.A2(g10512B),.A1(g4141B));
OR2_X1 U_g10558B (.ZN(g10558B),.A2(g10510B),.A1(g4126B));
OR2_X1 U_g11338B (.ZN(g11338B),.A2(g11178B),.A1(g11283B));
OR2_X1 U_g8435B (.ZN(g8435B),.A2(g8075B),.A1(g8403B));
OR2_X1 U_g10544B (.ZN(g10544B),.A2(g10495B),.A1(g4271B));
OR2_X1 U_g6911B (.ZN(g6911B),.A2(g5681B),.A1(g6342B));
OR2_X1 U_g10865B (.ZN(g10865B),.A2(g10752B),.A1(g5538B));
OR2_X1 U_g3698B (.ZN(g3698B),.A2(g869B),.A1(g3121B));
OR2_X1 U_g8214B (.ZN(g8214B),.A2(g7682B),.A1(g7472B));
OR2_X1 U_g6124B (.ZN(g6124B),.A2(g5188B),.A1(g5181B));
OR2_X1 U_g6469B (.ZN(g6469B),.A2(g4959B),.A1(g5698B));
OR2_X1 U_g5587B (.ZN(g5587B),.A2(g3904B),.A1(g4714B));
OR2_X1 U_g6177B (.ZN(g6177B),.A2(g4712B),.A1(g5444B));
OR2_X1 U_g9891B (.ZN(g9891B),.A2(g9760B),.A1(FE_OFN33_g9454B));
OR2_X1 U_g9913B (.ZN(g9913B),.A2(g9691B),.A1(g9849B));
OR4_X1 U_I5600B (.ZN(I5600B),.A4(g481B),.A3(g486B),.A2(g491B),.A1(g496B));
OR2_X1 U_g11257B (.ZN(g11257B),.A2(g11019B),.A1(g11234B));
OR2_X1 U_g8236B (.ZN(g8236B),.A2(g7680B),.A1(g7526B));
OR2_X1 U_g7385B (.ZN(g7385B),.A2(g6746B),.A1(g7235B));
OR2_X1 U_g6898B (.ZN(g6898B),.A2(g4881B),.A1(g6790B));
OR2_X1 U_g6900B (.ZN(g6900B),.A2(g6246B),.A1(g6787B));
OR2_X1 U_g4264B (.ZN(g4264B),.A2(g4053B),.A1(g4048B));
OR3_X1 U_g9726B (.ZN(g9726B),.A3(g9426B),.A2(g9420B),.A1(g9411B));
OR2_X1 U_g6088B (.ZN(g6088B),.A2(g4522B),.A1(g5260B));
OR2_X1 U_g6923B (.ZN(g6923B),.A2(g5695B),.A1(g6353B));
OR2_X1 U_g8194B (.ZN(g8194B),.A2(g7940B),.A1(g5168B));
OR3_X1 U_g9676B (.ZN(g9676B),.A3(FE_OFN62_g9274B),.A2(FE_OFN72_g9292B),.A1(g9454B));
OR2_X1 U_g11256B (.ZN(g11256B),.A2(g11018B),.A1(g11186B));
OR2_X1 U_g3860B (.ZN(g3860B),.A2(g2167B),.A1(g3107B));
OR2_X1 U_g11280B (.ZN(g11280B),.A2(g11153B),.A1(g11254B));
OR4_X1 U_g9727B (.ZN(g9727B),.A4(I14866B),.A3(g9391B),.A2(g9663B),.A1(g9650B));
OR2_X1 U_g4997B (.ZN(g4997B),.A2(g4584B),.A1(g4581B));
OR2_X1 U_g11624B (.ZN(g11624B),.A2(g11571B),.A1(g11595B));
OR2_X1 U_g11300B (.ZN(g11300B),.A2(g11091B),.A1(g11213B));
OR2_X1 U_g4238B (.ZN(g4238B),.A2(g4007B),.A1(g3999B));
OR2_X1 U_g8814B (.ZN(g8814B),.A2(g8728B),.A1(g7945B));
OR2_X1 U_g10401B (.ZN(g10401B),.A2(g10291B),.A1(g9317B));
OR2_X1 U_g8773B (.ZN(g8773B),.A2(g8653B),.A1(g5491B));
OR2_X1 U_g11231B (.ZN(g11231B),.A2(g11013B),.A1(g11156B));
OR2_X1 U_g10864B (.ZN(g10864B),.A2(g10751B),.A1(g5532B));
OR2_X1 U_g9624B (.ZN(g9624B),.A2(g9313B),.A1(g9316B));
OR3_X1 U_g9953B (.ZN(g9953B),.A3(g9803B),.A2(g9939B),.A1(g9945B));
OR2_X1 U_g6122B (.ZN(g6122B),.A2(g5180B),.A1(g5172B));
OR2_X1 U_g6465B (.ZN(g6465B),.A2(g5041B),.A1(g5825B));
OR2_X1 U_g6934B (.ZN(g6934B),.A2(g5720B),.A1(g6363B));
OR2_X1 U_g7664B (.ZN(g7664B),.A2(FE_OFN350_g3121B),.A1(g6855B));
OR2_X1 U_g7246B (.ZN(g7246B),.A2(g6003B),.A1(g6465B));
OR2_X1 U_g7203B (.ZN(g7203B),.A2(g6058B),.A1(g6640B));
OR2_X1 U_g6096B (.ZN(g6096B),.A2(g4542B),.A1(g5268B));
OR2_X1 U_g9747B (.ZN(g9747B),.A2(g9509B),.A1(g9173B));
OR2_X1 U_g11314B (.ZN(g11314B),.A2(g11102B),.A1(g11224B));
OR2_X1 U_g10733B (.ZN(g10733B),.A2(g10679B),.A1(g5227B));
OR2_X1 U_g8921B (.ZN(g8921B),.A2(g8748B),.A1(g8827B));
OR4_X1 U_I15054B (.ZN(I15054B),.A4(FE_OFN35_g9785B),.A3(FE_OFN61_g9624B),.A2(FE_OFN32_g9454B),.A1(FE_OFN90_I11360B));
OR2_X1 U_g11269B (.ZN(g11269B),.A2(g11031B),.A1(g11196B));
OR2_X1 U_g5555B (.ZN(g5555B),.A2(g4397B),.A1(g4389B));
OR2_X1 U_g11268B (.ZN(g11268B),.A2(g11030B),.A1(g11194B));
OR2_X1 U_g10485B (.ZN(g10485B),.A2(g10363B),.A1(g9317B));
OR2_X1 U_g10555B (.ZN(g10555B),.A2(g10504B),.A1(g4103B));
OR2_X1 U_g6481B (.ZN(g6481B),.A2(g4972B),.A1(g5722B));
OR2_X1 U_g10712B (.ZN(g10712B),.A2(g9097B),.A1(g10662B));
OR2_X1 U_g11335B (.ZN(g11335B),.A2(g11175B),.A1(g11279B));
OR2_X1 U_g8249B (.ZN(g8249B),.A2(g7710B),.A1(g8018B));
OR2_X1 U_g7638B (.ZN(g7638B),.A2(FE_OFN195_g6488B),.A1(g7265B));
OR2_X1 U_g10567B (.ZN(g10567B),.A2(g7378B),.A1(g10514B));
OR2_X1 U_g11487B (.ZN(g11487B),.A2(g11464B),.A1(g6662B));
OR4_X1 U_I15210B (.ZN(I15210B),.A4(g9882B),.A3(g9852B),.A2(g9964B),.A1(g9839B));
OR4_X1 U_I5805B (.ZN(I5805B),.A4(g2088B),.A3(g2096B),.A2(g2099B),.A1(g2102B));
OR2_X1 U_g8941B (.ZN(g8941B),.A2(FE_OFN332_g8748B),.A1(g8796B));
OR2_X1 U_g11443B (.ZN(g11443B),.A2(g11407B),.A1(g7130B));
OR2_X1 U_g4231B (.ZN(g4231B),.A2(g3998B),.A1(g3991B));
OR2_X1 U_g11278B (.ZN(g11278B),.A2(g11150B),.A1(g11253B));
OR2_X1 U_g11286B (.ZN(g11286B),.A2(g11209B),.A1(g10670B));
OR2_X1 U_g8431B (.ZN(g8431B),.A2(g8071B),.A1(g8387B));
OR2_X1 U_g7133B (.ZN(g7133B),.A2(I6273B),.A1(g6616B));
OR2_X1 U_g11306B (.ZN(g11306B),.A2(g11095B),.A1(g11216B));
OR2_X1 U_g8252B (.ZN(g8252B),.A2(g7679B),.A1(g7988B));
OR2_X1 U_g8812B (.ZN(g8812B),.A2(g8724B),.A1(g7939B));
OR2_X1 U_g7846B (.ZN(g7846B),.A2(g7241B),.A1(g7722B));
OR2_X1 U_g3875B (.ZN(g3875B),.A2(g12B),.A1(g3275B));
OR2_X1 U_g5996B (.ZN(g5996B),.A2(g3383B),.A1(g5473B));
OR2_X1 U_g6592B (.ZN(g6592B),.A2(g5882B),.A1(g5100B));
OR2_X1 U_g8286B (.ZN(g8286B),.A2(g7823B),.A1(g8107B));
OR2_X1 U_g10501B (.ZN(g10501B),.A2(g10445B),.A1(g4161B));
OR2_X1 U_g10728B (.ZN(g10728B),.A2(g10642B),.A1(g4973B));
OR2_X1 U_g8270B (.ZN(g8270B),.A2(g3434B),.A1(g7894B));
OR2_X1 U_g7290B (.ZN(g7290B),.A2(g6316B),.A1(g7046B));
OR2_X1 U_g6068B (.ZN(g6068B),.A2(g4497B),.A1(g5220B));
OR2_X1 U_g6468B (.ZN(g6468B),.A2(g4950B),.A1(g5690B));
OR2_X1 U_g11217B (.ZN(g11217B),.A2(g11005B),.A1(g11144B));
OR2_X1 U_g11478B (.ZN(g11478B),.A2(g11455B),.A1(g6532B));
OR4_X2 U_g9536B (.ZN(g9536B),.A4(g9324B),.A3(g9328B),.A2(g9331B),.A1(g9335B));
OR2_X1 U_g5981B (.ZN(g5981B),.A2(g4383B),.A1(g5074B));
OR2_X1 U_g11486B (.ZN(g11486B),.A2(g11463B),.A1(g6654B));
OR2_X1 U_g8377B (.ZN(g8377B),.A2(g7958B),.A1(g8185B));
OR2_X1 U_g8206B (.ZN(g8206B),.A2(g7683B),.A1(g7459B));
OR2_X1 U_g11580B (.ZN(g11580B),.A2(g11544B),.A1(g11413B));
OR2_X1 U_g8287B (.ZN(g8287B),.A2(g7824B),.A1(g8117B));
OR2_X1 U_g11223B (.ZN(g11223B),.A2(g11008B),.A1(g11147B));
OR2_X1 U_g9522B (.ZN(g9522B),.A2(FE_OFN44_g9125B),.A1(g9173B));
OR2_X1 U_g8199B (.ZN(g8199B),.A2(g7444B),.A1(g7902B));
OR2_X1 U_g5802B (.ZN(g5802B),.A2(g4837B),.A1(g5601B));
OR2_X1 U_g11321B (.ZN(g11321B),.A2(g11105B),.A1(g11230B));
OR2_X1 U_g6524B (.ZN(g6524B),.A2(g4996B),.A1(g5746B));
OR2_X1 U_g10664B (.ZN(g10664B),.A2(g10582B),.A1(g10240B));
OR2_X1 U_g7257B (.ZN(g7257B),.A2(g4725B),.A1(g6701B));
OR2_X1 U_g7301B (.ZN(g7301B),.A2(g6327B),.A1(g7140B));
OR2_X1 U_g10484B (.ZN(g10484B),.A2(g10400B),.A1(g9317B));
OR2_X1 U_g10554B (.ZN(g10554B),.A2(g10503B),.A1(g4097B));
OR2_X1 U_g8259B (.ZN(g8259B),.A2(g7719B),.A1(g8028B));
OR2_X1 U_g11334B (.ZN(g11334B),.A2(g11174B),.A1(g11277B));
OR2_X1 U_g8819B (.ZN(g8819B),.A2(g8734B),.A1(g7957B));
OR2_X1 U_g8923B (.ZN(g8923B),.A2(FE_OFN329_g8763B),.A1(g8846B));
OR2_X2 U_g8488B (.ZN(g8488B),.A2(g8390B),.A1(FE_OFN204_g3664B));
OR2_X1 U_g7441B (.ZN(g7441B),.A2(g5867B),.A1(g7271B));
OR2_X1 U_g6026B (.ZN(g6026B),.A2(g3970B),.A1(g5507B));
OR2_X1 U_g10799B (.ZN(g10799B),.A2(g10769B),.A1(g6225B));
OR2_X1 U_g10798B (.ZN(g10798B),.A2(g10768B),.A1(g6217B));
OR2_X1 U_g10805B (.ZN(g10805B),.A2(g10760B),.A1(g10759B));
OR2_X1 U_g10732B (.ZN(g10732B),.A2(g10661B),.A1(g4358B));
OR2_X1 U_g6061B (.ZN(g6061B),.A2(g4B),.A1(g5204B));
OR2_X1 U_g9512B (.ZN(g9512B),.A2(g9125B),.A1(g9151B));
OR2_X1 U_g10013B (.ZN(g10013B),.A2(I15215B),.A1(I15214B));
OR2_X1 U_g8806B (.ZN(g8806B),.A2(g8718B),.A1(g7931B));
OR2_X1 U_g8943B (.ZN(g8943B),.A2(FE_OFN332_g8748B),.A1(g8837B));
OR2_X1 U_g11293B (.ZN(g11293B),.A2(g10818B),.A1(g11211B));
OR2_X1 U_g11265B (.ZN(g11265B),.A2(g11027B),.A1(g11189B));
OR2_X1 U_g8887B (.ZN(g8887B),.A2(FE_OFN329_g8763B),.A1(g8842B));
OR2_X1 U_g5838B (.ZN(g5838B),.A2(g3974B),.A1(g5612B));
OR2_X1 U_g6514B (.ZN(g6514B),.A2(g4992B),.A1(g5738B));
OR2_X1 U_g8322B (.ZN(g8322B),.A2(g6891B),.A1(g8136B));
OR2_X1 U_g8230B (.ZN(g8230B),.A2(g7686B),.A1(g7515B));
OR2_X1 U_g5809B (.ZN(g5809B),.A2(g4865B),.A1(g5611B));
OR2_X1 U_g8433B (.ZN(g8433B),.A2(g8073B),.A1(g8399B));
OR2_X1 U_g11579B (.ZN(g11579B),.A2(g11551B),.A1(g5123B));
OR2_X1 U_g10771B (.ZN(g10771B),.A2(g10684B),.A1(g5533B));
OR2_X1 U_g11615B (.ZN(g11615B),.A2(g11592B),.A1(g11601B));
OR2_X1 U_g9367B (.ZN(g9367B),.A2(g9331B),.A1(g9335B));
OR3_X1 U_g9872B (.ZN(g9872B),.A3(g9759B),.A2(g9594B),.A1(g9617B));
OR2_X1 U_g6522B (.ZN(g6522B),.A2(g4994B),.A1(g5744B));
OR2_X1 U_g8266B (.ZN(g8266B),.A2(g3412B),.A1(g7885B));
OR2_X1 U_g10414B (.ZN(g10414B),.A2(g9291B),.A1(g10300B));
OR2_X1 U_g11275B (.ZN(g11275B),.A2(g11148B),.A1(g11248B));
OR2_X1 U_g11430B (.ZN(g11430B),.A2(g4006B),.A1(g11387B));
OR2_X1 U_g8248B (.ZN(g8248B),.A2(g7707B),.A1(g8014B));
OR2_X1 U_g8815B (.ZN(g8815B),.A2(g8730B),.A1(g7948B));
OR2_X1 U_g7183B (.ZN(g7183B),.A2(I9717B),.A1(g6623B));
OR2_X1 U_g5983B (.ZN(g5983B),.A2(g4392B),.A1(g5084B));
OR2_X1 U_g8154B (.ZN(g8154B),.A2(g6879B),.A1(g7891B));
OR2_X1 U_g6537B (.ZN(g6537B),.A2(g5005B),.A1(g5781B));
OR2_X1 U_g4309B (.ZN(g4309B),.A2(g4079B),.A1(g4069B));
OR2_X1 U_g10725B (.ZN(g10725B),.A2(g10634B),.A1(g4962B));
OR2_X1 U_g6243B (.ZN(g6243B),.A2(g4144B),.A1(g5537B));
OR4_X1 U_I6351B (.ZN(I6351B),.A4(g2372B),.A3(g2380B),.A2(g2389B),.A1(g2405B));
OR3_X1 U_g9519B (.ZN(g9519B),.A3(FE_OFN44_g9125B),.A2(g9151B),.A1(g9173B));
OR2_X1 U_g9740B (.ZN(g9740B),.A2(g9505B),.A1(g9418B));
OR2_X1 U_g8267B (.ZN(g8267B),.A2(g3422B),.A1(g7889B));
OR3_X1 U_g10744B (.ZN(g10744B),.A3(I16427B),.A2(g10668B),.A1(g10381B));
OR2_X1 U_g6542B (.ZN(g6542B),.A2(g5010B),.A1(g5789B));
OR2_X1 U_g7303B (.ZN(g7303B),.A2(g6329B),.A1(g7145B));
OR2_X1 U_g10652B (.ZN(g10652B),.A2(g7743B),.A1(g10627B));
OR2_X1 U_g5036B (.ZN(g5036B),.A2(g4162B),.A1(g4871B));
OR2_X1 U_g7240B (.ZN(g7240B),.A2(g6095B),.A1(g6687B));
OR2_X1 U_g8221B (.ZN(g8221B),.A2(g7688B),.A1(g7496B));
OR2_X1 U_g6902B (.ZN(g6902B),.A2(g4223B),.A1(g6794B));
OR2_X1 U_g10500B (.ZN(g10500B),.A2(g10442B),.A1(g4157B));
OR2_X1 U_g4052B (.ZN(g4052B),.A2(g2515B),.A1(g2862B));
OR4_X1 U_I14858B (.ZN(I14858B),.A4(g9602B),.A3(g9610B),.A2(g9595B),.A1(g9585B));
OR2_X1 U_g6529B (.ZN(g6529B),.A2(g5000B),.A1(g5757B));
OR2_X1 U_g11264B (.ZN(g11264B),.A2(g11026B),.A1(g11188B));
OR4_X1 U_I15209B (.ZN(I15209B),.A4(g9830B),.A3(g9934B),.A2(g9905B),.A1(g8169B));
OR2_X1 U_g8241B (.ZN(g8241B),.A2(g7684B),.A1(g7536B));
OR2_X1 U_g10795B (.ZN(g10795B),.A2(g10764B),.A1(g6199B));
OR2_X1 U_g11607B (.ZN(g11607B),.A2(g11557B),.A1(g11586B));
OR2_X1 U_g8644B (.ZN(g8644B),.A2(g8464B),.A1(g8123B));
OR3_X1 U_g4682B (.ZN(g4682B),.A3(g1570B),.A2(g3348B),.A1(g3563B));
OR2_X1 U_g8818B (.ZN(g8818B),.A2(g8733B),.A1(g7955B));
OR2_X1 U_g2984B (.ZN(g2984B),.A2(g2522B),.A1(g2528B));
OR2_X1 U_g9931B (.ZN(g9931B),.A2(g9900B),.A1(g8931B));
OR2_X1 U_g3414B (.ZN(g3414B),.A2(g2917B),.A1(g2911B));
OR2_X1 U_g9515B (.ZN(g9515B),.A2(g9151B),.A1(g9173B));
OR2_X1 U_g10724B (.ZN(g10724B),.A2(g10672B),.A1(g10312B));
OR2_X1 U_g7294B (.ZN(g7294B),.A2(g6320B),.A1(g7068B));
OR2_X1 U_g5189B (.ZN(g5189B),.A2(FE_OFN292_g3015B),.A1(g4345B));
OR2_X1 U_g8614B (.ZN(g8614B),.A2(g8510B),.A1(g8365B));
OR2_X1 U_g3513B (.ZN(g3513B),.A2(g2180B),.A1(g3118B));
OR2_X1 U_g6909B (.ZN(g6909B),.A2(g5309B),.A1(g6346B));
OR4_X1 U_I5571B (.ZN(I5571B),.A4(g426B),.A3(g386B),.A2(g391B),.A1(g396B));
OR2_X1 U_g4283B (.ZN(g4283B),.A2(g4063B),.A1(g4059B));
OR2_X1 U_g8939B (.ZN(g8939B),.A2(FE_OFN332_g8748B),.A1(g8791B));
OR2_X1 U_g2514B (.ZN(g2514B),.A2(I5600B),.A1(I5599B));
OR2_X1 U_g11327B (.ZN(g11327B),.A2(g11167B),.A1(g11297B));
OR2_X1 U_g8187B (.ZN(g8187B),.A2(g7677B),.A1(g7542B));
OR2_X1 U_g11606B (.ZN(g11606B),.A2(g11556B),.A1(g11585B));
OR2_X1 U_g11303B (.ZN(g11303B),.A2(g11092B),.A1(g11214B));
OR2_X1 U_g5309B (.ZN(g5309B),.A2(g4401B),.A1(FE_OFN204_g3664B));
OR2_X1 U_g8200B (.ZN(g8200B),.A2(g7685B),.A1(g7535B));
OR3_X1 U_g2522B (.ZN(g2522B),.A3(I5629B),.A2(g829B),.A1(g833B));
OR4_X1 U_g2315B (.ZN(g2315B),.A4(I5363B),.A3(g1113B),.A2(g1166B),.A1(g1163B));
OR2_X1 U_g6506B (.ZN(g6506B),.A2(g4989B),.A1(g5731B));
OR2_X1 U_g10649B (.ZN(g10649B),.A2(g7741B),.A1(g10626B));
OR2_X1 U_g8159B (.ZN(g8159B),.A2(g6886B),.A1(g7895B));
OR2_X1 U_g7626B (.ZN(g7626B),.A2(g3440B),.A1(g7060B));
OR2_X1 U_g10770B (.ZN(g10770B),.A2(g10682B),.A1(g5525B));
OR2_X1 U_g11483B (.ZN(g11483B),.A2(g11460B),.A1(g6633B));
OR2_X1 U_g8811B (.ZN(g8811B),.A2(g8722B),.A1(g7935B));
OR3_X1 U_g8642B (.ZN(g8642B),.A3(g8465B),.A2(g31B),.A1(g30B));
OR2_X1 U_g6545B (.ZN(g6545B),.A2(g5025B),.A1(g5795B));
OR2_X1 U_g10767B (.ZN(g10767B),.A2(g10681B),.A1(g5500B));
OR2_X1 U_g11326B (.ZN(g11326B),.A2(g11166B),.A1(g11296B));
OR2_X1 U_g10898B (.ZN(g10898B),.A2(g10777B),.A1(g4220B));
OR2_X1 U_g11252B (.ZN(g11252B),.A2(g10969B),.A1(g11099B));
OR2_X1 U_g10719B (.ZN(g10719B),.A2(g10666B),.A1(g10303B));
OR2_X1 U_g4609B (.ZN(g4609B),.A2(g119B),.A1(g3275B));
OR2_X1 U_g6507B (.ZN(g6507B),.A2(g4990B),.A1(g5732B));
OR2_X1 U_g10718B (.ZN(g10718B),.A2(g10706B),.A1(g6238B));
OR2_X1 U_g10521B (.ZN(g10521B),.A2(I16149B),.A1(I16148B));
OR2_X1 U_g7075B (.ZN(g7075B),.A2(g6530B),.A1(g5104B));
OR2_X1 U_g7292B (.ZN(g7292B),.A2(g6318B),.A1(g7055B));
OR2_X1 U_g10861B (.ZN(g10861B),.A2(g10745B),.A1(g5523B));
OR2_X1 U_g8417B (.ZN(g8417B),.A2(g7721B),.A1(g8246B));
OR2_X1 U_g6515B (.ZN(g6515B),.A2(g4993B),.A1(g5739B));
OR4_X1 U_I14855B (.ZN(I14855B),.A4(g9596B),.A3(g9601B),.A2(g9593B),.A1(g9583B));
OR4_X1 U_I15205B (.ZN(I15205B),.A4(g9878B),.A3(g9850B),.A2(g9963B),.A1(g9838B));
OR4_X1 U_I15051B (.ZN(I15051B),.A4(FE_OFN35_g9785B),.A3(FE_OFN60_g9624B),.A2(g9673B),.A1(FE_OFN90_I11360B));
OR3_X1 U_g9724B (.ZN(g9724B),.A3(g9426B),.A2(g9419B),.A1(g9409B));
OR2_X1 U_g6528B (.ZN(g6528B),.A2(g4999B),.A1(g5756B));
OR2_X1 U_g8823B (.ZN(g8823B),.A2(g8693B),.A1(g8778B));
OR2_X1 U_g7503B (.ZN(g7503B),.A2(g6430B),.A1(g6887B));
OR2_X1 U_g8148B (.ZN(g8148B),.A2(g6872B),.A1(g7884B));
OR2_X1 U_g8649B (.ZN(g8649B),.A2(g3440B),.A1(g8499B));
OR2_X1 U_g3584B (.ZN(g3584B),.A2(g2516B),.A1(g2863B));
OR2_X1 U_g10776B (.ZN(g10776B),.A2(g10758B),.A1(g5544B));
OR3_X1 U_g9680B (.ZN(g9680B),.A3(FE_OFN62_g9274B),.A2(FE_OFN72_g9292B),.A1(FE_OFN32_g9454B));
OR2_X1 U_g10859B (.ZN(g10859B),.A2(g10742B),.A1(g5512B));
OR3_X1 U_I14866B (.ZN(I14866B),.A3(g9619B),.A2(g9609B),.A1(g9590B));
OR2_X1 U_g7299B (.ZN(g7299B),.A2(g6325B),.A1(g7138B));
OR2_X1 U_g10858B (.ZN(g10858B),.A2(g10741B),.A1(g5501B));
OR2_X1 U_g8193B (.ZN(g8193B),.A2(g7937B),.A1(g5145B));
OR3_X1 U_g9511B (.ZN(g9511B),.A3(g9111B),.A2(g9125B),.A1(g9151B));
OR2_X1 U_g7738B (.ZN(g7738B),.A2(g6738B),.A1(g7200B));
OR2_X1 U_g7244B (.ZN(g7244B),.A2(g4720B),.A1(g6699B));
OR2_X1 U_g3425B (.ZN(g3425B),.A2(g2910B),.A1(g2895B));
OR2_X1 U_g7478B (.ZN(g7478B),.A2(g6423B),.A1(g6884B));
OR3_X1 U_g9714B (.ZN(g9714B),.A3(g9654B),.A2(g9366B),.A1(g9664B));
OR2_X1 U_g10025B (.ZN(g10025B),.A2(I15225B),.A1(I15224B));
OR2_X1 U_g6908B (.ZN(g6908B),.A2(g4229B),.A1(g6345B));
OR2_X1 U_g5028B (.ZN(g5028B),.A2(g4128B),.A1(g4836B));
OR2_X1 U_g8253B (.ZN(g8253B),.A2(g7718B),.A1(g8023B));
OR2_X1 U_g8938B (.ZN(g8938B),.A2(FE_OFN332_g8748B),.A1(g8789B));
OR2_X1 U_g8813B (.ZN(g8813B),.A2(g8726B),.A1(g7943B));
OR2_X1 U_g9736B (.ZN(g9736B),.A2(g9423B),.A1(g9430B));
OR2_X1 U_g9968B (.ZN(g9968B),.A2(I15172B),.A1(I15171B));
OR2_X1 U_g8552B (.ZN(g8552B),.A2(g8388B),.A1(g8217B));
OR2_X1 U_g5910B (.ZN(g5910B),.A2(g4341B),.A1(g5023B));
OR2_X1 U_g11249B (.ZN(g11249B),.A2(g11143B),.A1(g6162B));
OR2_X1 U_g11482B (.ZN(g11482B),.A2(g11459B),.A1(g6628B));
OR4_X1 U_g9722B (.ZN(g9722B),.A4(I14855B),.A3(g9391B),.A2(g9643B),.A1(g9612B));
OR4_X1 U_I15204B (.ZN(I15204B),.A4(g9829B),.A3(g9933B),.A2(g9904B),.A1(g8168B));
OR2_X1 U_g7236B (.ZN(g7236B),.A2(g6092B),.A1(g6684B));
OR2_X1 U_g8645B (.ZN(g8645B),.A2(g8469B),.A1(g8127B));
OR2_X1 U_g11647B (.ZN(g11647B),.A2(g11637B),.A1(g6622B));
OR2_X1 U_g6777B (.ZN(g6777B),.A2(g48B),.A1(I9221B));
OR3_X1 U_g9737B (.ZN(g9737B),.A3(g9387B),.A2(g9658B),.A1(g9657B));
OR4_X1 U_I16149B (.ZN(I16149B),.A4(g10467B),.A3(g10468B),.A2(g10470B),.A1(g10472B));
OR2_X1 U_g11233B (.ZN(g11233B),.A2(g10946B),.A1(g11085B));
OR2_X1 U_g8607B (.ZN(g8607B),.A2(g8554B),.A1(g8406B));
OR4_X1 U_I16148B (.ZN(I16148B),.A4(g10474B),.A3(g10476B),.A2(g10384B),.A1(g10386B));
OR2_X1 U_g8158B (.ZN(g8158B),.A2(g6883B),.A1(g7893B));
OR2_X1 U_g5846B (.ZN(g5846B),.A2(g4236B),.A1(g4932B));
OR2_X1 U_g5396B (.ZN(g5396B),.A2(g3684B),.A1(g4481B));
OR2_X1 U_g5803B (.ZN(g5803B),.A2(g3383B),.A1(g5575B));
OR2_X1 U_g11331B (.ZN(g11331B),.A2(g11171B),.A1(g11272B));
OR2_X1 U_g7295B (.ZN(g7295B),.A2(g6321B),.A1(g7071B));
OR2_X1 U_g6541B (.ZN(g6541B),.A2(g5009B),.A1(g5788B));
OR2_X1 U_g8615B (.ZN(g8615B),.A2(g8557B),.A1(g8413B));
OR2_X1 U_g9926B (.ZN(g9926B),.A2(g9715B),.A1(g9868B));
OR2_X1 U_g9754B (.ZN(g9754B),.A2(g9511B),.A1(g9173B));
OR2_X1 U_g8284B (.ZN(g8284B),.A2(g7821B),.A1(g8102B));
OR2_X1 U_g2204B (.ZN(g2204B),.A2(g1394B),.A1(g1393B));
OR2_X1 U_g7471B (.ZN(g7471B),.A2(g6416B),.A1(g6880B));
OR2_X1 U_g7242B (.ZN(g7242B),.A2(g6098B),.A1(g6693B));
OR2_X1 U_g5847B (.ZN(g5847B),.A2(g3987B),.A1(g5626B));
OR2_X1 U_g6901B (.ZN(g6901B),.A2(g6247B),.A1(g6788B));
OR2_X1 U_g8559B (.ZN(g8559B),.A2(g3664B),.A1(g8380B));
OR3_X1 U_g9729B (.ZN(g9729B),.A3(g9387B),.A2(g9357B),.A1(g9618B));
OR2_X1 U_g10860B (.ZN(g10860B),.A2(g10743B),.A1(g5513B));
OR2_X1 U_g9927B (.ZN(g9927B),.A2(g9716B),.A1(g9869B));
OR2_X1 U_g10497B (.ZN(g10497B),.A2(g10396B),.A1(FE_OFN277_g48B));
OR4_X1 U_g9885B (.ZN(g9885B),.A4(g9759B),.A3(g9662B),.A2(g9598B),.A1(g9454B));
OR4_X1 U_g2528B (.ZN(g2528B),.A4(g849B),.A3(g853B),.A2(g857B),.A1(g861B));
OR2_X1 U_g11229B (.ZN(g11229B),.A2(g11012B),.A1(g11154B));
OR2_X1 U_g8973B (.ZN(g8973B),.A2(FE_OFN329_g8763B),.A1(g8821B));
OR2_X1 U_g10658B (.ZN(g10658B),.A2(g7674B),.A1(g10595B));
OR2_X1 U_g10339B (.ZN(g10339B),.A2(g9291B),.A1(g10232B));
OR4_X1 U_I5363B (.ZN(I5363B),.A4(g1160B),.A3(g1157B),.A2(g1153B),.A1(g1149B));
OR2_X1 U_g11310B (.ZN(g11310B),.A2(g11100B),.A1(g11220B));
OR2_X1 U_g6500B (.ZN(g6500B),.A2(g4986B),.A1(g5725B));
OR2_X1 U_g10855B (.ZN(g10855B),.A2(g10736B),.A1(g6075B));
OR2_X1 U_g9916B (.ZN(g9916B),.A2(g9694B),.A1(g9855B));
OR2_X1 U_g10411B (.ZN(g10411B),.A2(g9291B),.A1(g10299B));
OR2_X1 U_g11603B (.ZN(g11603B),.A2(g11553B),.A1(g11582B));
OR4_X1 U_I5357B (.ZN(I5357B),.A4(g1250B),.A3(g1255B),.A2(g1260B),.A1(g1265B));
OR2_X1 U_g6672B (.ZN(g6672B),.A2(g5259B),.A1(g5509B));
OR3_X1 U_g9873B (.ZN(g9873B),.A3(g9758B),.A2(g9599B),.A1(g9623B));
OR2_X1 U_g6523B (.ZN(g6523B),.A2(g4995B),.A1(g5745B));
OR2_X1 U_g10707B (.ZN(g10707B),.A2(g10686B),.A1(g5545B));
OR4_X1 U_I5626B (.ZN(I5626B),.A4(g534B),.A3(g530B),.A2(g525B),.A1(g521B));
OR2_X1 U_g9579B (.ZN(g9579B),.A2(g9030B),.A1(FE_OFN54_g9052B));
OR2_X1 U_g7298B (.ZN(g7298B),.A2(g6324B),.A1(g7136B));
OR2_X1 U_g6551B (.ZN(g6551B),.A2(g5031B),.A1(g5804B));
OR2_X1 U_g6099B (.ZN(g6099B),.A2(g4550B),.A1(g5273B));
OR2_X1 U_g8282B (.ZN(g8282B),.A2(g7819B),.A1(g8101B));
OR2_X1 U_g9917B (.ZN(g9917B),.A2(g9695B),.A1(g9856B));
OR4_X1 U_I15057B (.ZN(I15057B),.A4(FE_OFN35_g9785B),.A3(FE_OFN60_g9624B),.A2(g9680B),.A1(FE_OFN90_I11360B));
OR2_X1 U_g7219B (.ZN(g7219B),.A2(I9717B),.A1(g6661B));
OR2_X1 U_g10019B (.ZN(g10019B),.A2(I15220B),.A1(I15219B));
OR2_X1 U_g5857B (.ZN(g5857B),.A2(g4670B),.A1(g5418B));
OR4_X1 U_g9725B (.ZN(g9725B),.A4(I14862B),.A3(g9391B),.A2(g9659B),.A1(g9642B));
OR2_X1 U_g11298B (.ZN(g11298B),.A2(g11087B),.A1(g11212B));
OR2_X1 U_g10402B (.ZN(g10402B),.A2(g9291B),.A1(g10295B));
OR4_X1 U_g2521B (.ZN(g2521B),.A4(I5626B),.A3(g476B),.A2(g542B),.A1(g538B));
OR2_X1 U_g10866B (.ZN(g10866B),.A2(g10753B),.A1(g5539B));
OR2_X1 U_g6534B (.ZN(g6534B),.A2(g5003B),.A1(g5772B));
OR2_X1 U_g11232B (.ZN(g11232B),.A2(g11015B),.A1(g11158B));
OR3_X1 U_g9706B (.ZN(g9706B),.A3(g9591B),.A2(g9386B),.A1(g9644B));
OR2_X1 U_g10001B (.ZN(g10001B),.A2(I15205B),.A1(I15204B));
OR2_X1 U_g8776B (.ZN(g8776B),.A2(g8655B),.A1(g5510B));
OR2_X1 U_g7225B (.ZN(g7225B),.A2(g6079B),.A1(g6666B));
OR3_X1 U_g9888B (.ZN(g9888B),.A3(g9757B),.A2(g9608B),.A1(g9648B));
OR2_X1 U_g11261B (.ZN(g11261B),.A2(g11023B),.A1(g11238B));
OR3_X1 U_g9956B (.ZN(g9956B),.A3(g9815B),.A2(g9942B),.A1(g9948B));
OR2_X1 U_g10923B (.ZN(g10923B),.A2(g10715B),.A1(g10778B));
OR2_X1 U_g8264B (.ZN(g8264B),.A2(g3912B),.A1(g7879B));
OR2_X1 U_g6513B (.ZN(g6513B),.A2(g4991B),.A1(g5737B));
OR3_X1 U_I14835B (.ZN(I14835B),.A3(g9588B),.A2(g9645B),.A1(g9621B));
OR2_X1 U_g8641B (.ZN(g8641B),.A2(g8463B),.A1(g8120B));
OR3_X1 U_g5361B (.ZN(g5361B),.A3(g126B),.A2(g3348B),.A1(g4316B));
OR2_X1 U_g11316B (.ZN(g11316B),.A2(g11103B),.A1(g11226B));
OR4_X1 U_I16161B (.ZN(I16161B),.A4(g10475B),.A3(g10477B),.A2(g10478B),.A1(g10479B));
OR2_X1 U_g6916B (.ZN(g6916B),.A2(g5687B),.A1(g6348B));
OR2_X1 U_g8777B (.ZN(g8777B),.A2(g8659B),.A1(g5522B));
OR4_X1 U_g2353B (.ZN(g2353B),.A4(g1415B),.A3(g1411B),.A2(g1407B),.A1(g1403B));
OR2_X1 U_g7510B (.ZN(g7510B),.A2(g6730B),.A1(g7186B));
OR3_X1 U_g9957B (.ZN(g9957B),.A3(g9803B),.A2(g9943B),.A1(g9949B));
OR2_X1 U_g2744B (.ZN(g2744B),.A2(I5805B),.A1(I5804B));
OR2_X1 U_g7245B (.ZN(g7245B),.A2(g6102B),.A1(g6696B));
OR2_X1 U_g7291B (.ZN(g7291B),.A2(g6317B),.A1(g7050B));
OR2_X1 U_g8611B (.ZN(g8611B),.A2(g8556B),.A1(g8410B));
OR4_X1 U_I15199B (.ZN(I15199B),.A4(g9828B),.A3(g9932B),.A2(g9903B),.A1(g8167B));
OR2_X1 U_g10550B (.ZN(g10550B),.A2(g10450B),.A1(g4437B));
OR2_X1 U_g11330B (.ZN(g11330B),.A2(g11170B),.A1(g11304B));
OR2_X1 U_g10721B (.ZN(g10721B),.A2(g10669B),.A1(g10306B));
OR2_X1 U_g8153B (.ZN(g8153B),.A2(g6875B),.A1(g7888B));
OR2_X1 U_g10773B (.ZN(g10773B),.A2(g10685B),.A1(g5540B));
OR2_X1 U_g3688B (.ZN(g3688B),.A2(g868B),.A1(g3744B));
OR4_X1 U_I15225B (.ZN(I15225B),.A4(g9881B),.A3(g9859B),.A2(g9967B),.A1(g9842B));
OR2_X1 U_g6042B (.ZN(g6042B),.A2(g3987B),.A1(g5535B));
OR2_X1 U_g10655B (.ZN(g10655B),.A2(g7389B),.A1(g10561B));
OR2_X1 U_g11259B (.ZN(g11259B),.A2(g11021B),.A1(g11236B));
OR2_X1 U_g11225B (.ZN(g11225B),.A2(g11009B),.A1(g11149B));
OR2_X1 U_g5914B (.ZN(g5914B),.A2(g4343B),.A1(g5029B));
OR2_X1 U_g11258B (.ZN(g11258B),.A2(g11020B),.A1(g11235B));
OR2_X1 U_g6054B (.ZN(g6054B),.A2(g4483B),.A1(g5199B));
OR3_X1 U_g9728B (.ZN(g9728B),.A3(g9426B),.A2(g9422B),.A1(g9412B));
OR3_X1 U_g9730B (.ZN(g9730B),.A3(g9423B),.A2(g9425B),.A1(g9414B));
OR2_X1 U_g5820B (.ZN(g5820B),.A2(g3942B),.A1(g5595B));
OR3_X1 U_g8574B (.ZN(g8574B),.A3(g8465B),.A2(I11360B),.A1(g30B));
OR2_X1 U_g11602B (.ZN(g11602B),.A2(g11552B),.A1(g11581B));
OR2_X1 U_g10502B (.ZN(g10502B),.A2(g10503B),.A1(g4169B));
OR2_X1 U_g10557B (.ZN(g10557B),.A2(g10508B),.A1(g4123B));
OR4_X1 U_I15171B (.ZN(I15171B),.A4(g9835B),.A3(g9896B),.A2(g9909B),.A1(g8175B));
OR2_X1 U_g11337B (.ZN(g11337B),.A2(g11177B),.A1(g11282B));
OR2_X1 U_g7465B (.ZN(g7465B),.A2(g6410B),.A1(g6876B));
OR2_X1 U_g8262B (.ZN(g8262B),.A2(g7625B),.A1(g7970B));
OR2_X1 U_g8889B (.ZN(g8889B),.A2(FE_OFN329_g8763B),.A1(g8844B));
OR2_X1 U_g7096B (.ZN(g7096B),.A2(g5911B),.A1(g6544B));
OR2_X1 U_g5995B (.ZN(g5995B),.A2(g5099B),.A1(g5097B));
OR2_X1 U_g8285B (.ZN(g8285B),.A2(g7822B),.A1(g8104B));
OR2_X1 U_g10791B (.ZN(g10791B),.A2(g10762B),.A1(g6186B));
OR2_X1 U_g2499B (.ZN(g2499B),.A2(I5571B),.A1(I5570B));
OR2_X1 U_g6049B (.ZN(g6049B),.A2(g4670B),.A1(g5254B));
OR2_X1 U_g9920B (.ZN(g9920B),.A2(g9701B),.A1(g9860B));
OR2_X1 U_g10556B (.ZN(g10556B),.A2(g10506B),.A1(g4115B));
OR2_X1 U_g8643B (.ZN(g8643B),.A2(g8508B),.A1(g8364B));
OR2_X1 U_g5810B (.ZN(g5810B),.A2(g3912B),.A1(g5588B));
OR2_X1 U_g11336B (.ZN(g11336B),.A2(g11176B),.A1(g11281B));
OR2_X1 U_g8742B (.ZN(g8742B),.A2(g8598B),.A1(g8135B));
OR2_X1 U_g8926B (.ZN(g8926B),.A2(g8763B),.A1(g8848B));
OR2_X1 U_g7218B (.ZN(g7218B),.A2(g6070B),.A1(g6655B));
OR4_X1 U_I15224B (.ZN(I15224B),.A4(g9834B),.A3(g9937B),.A2(g9908B),.A1(g8174B));
OR2_X1 U_g7293B (.ZN(g7293B),.A2(g6319B),.A1(g7063B));
OR2_X1 U_g11288B (.ZN(g11288B),.A2(g11070B),.A1(g11204B));
OR2_X1 U_g10800B (.ZN(g10800B),.A2(g10772B),.A1(g6245B));
OR2_X1 U_g11308B (.ZN(g11308B),.A2(g11098B),.A1(g11218B));
OR2_X1 U_g8269B (.ZN(g8269B),.A2(g3429B),.A1(g7892B));
OR2_X1 U_g10417B (.ZN(g10417B),.A2(g9097B),.A1(g10301B));
OR2_X1 U_g10936B (.ZN(g10936B),.A2(g10808B),.A1(g5170B));
OR2_X1 U_g9388B (.ZN(g9388B),.A2(g9223B),.A1(g9240B));
OR2_X1 U_g6185B (.ZN(g6185B),.A2(g4715B),.A1(g5470B));
OR2_X1 U_g6470B (.ZN(g6470B),.A2(g4960B),.A1(g5699B));
OR2_X1 U_g6897B (.ZN(g6897B),.A2(g6240B),.A1(g6771B));
OR2_X1 U_g8885B (.ZN(g8885B),.A2(FE_OFN329_g8763B),.A1(g8841B));
OR2_X1 U_g11260B (.ZN(g11260B),.A2(g11022B),.A1(g11237B));
OR2_X1 U_g11488B (.ZN(g11488B),.A2(g11465B),.A1(g6671B));
OR2_X1 U_g6105B (.ZN(g6105B),.A2(g4559B),.A1(g5279B));
OR2_X1 U_g10807B (.ZN(g10807B),.A2(g10761B),.A1(g10701B));
OR2_X1 U_g10639B (.ZN(g10639B),.A2(g7734B),.A1(g10623B));
OR2_X1 U_g4556B (.ZN(g4556B),.A2(g1212B),.A1(g3536B));
OR2_X1 U_g8288B (.ZN(g8288B),.A2(g7825B),.A1(g8119B));
OR2_X1 U_g6755B (.ZN(g6755B),.A2(g5479B),.A1(g4934B));
OR3_X1 U_I14862B (.ZN(I14862B),.A3(g9611B),.A2(g9600B),.A1(g9587B));
OR4_X1 U_I16160B (.ZN(I16160B),.A4(g10481B),.A3(g10482B),.A2(g10392B),.A1(g10394B));
OR2_X1 U_g11610B (.ZN(g11610B),.A2(g11560B),.A1(g11589B));
OR4_X1 U_g9711B (.ZN(g9711B),.A4(g9589B),.A3(g9359B),.A2(g9390B),.A1(g9660B));
OR2_X1 U_g6045B (.ZN(g6045B),.A2(g3989B),.A1(g5541B));
OR2_X1 U_g11270B (.ZN(g11270B),.A2(g11032B),.A1(g11198B));
OR2_X1 U_g7258B (.ZN(g7258B),.A2(g5913B),.A1(g6549B));
OR2_X1 U_g6059B (.ZN(g6059B),.A2(g4489B),.A1(g5211B));
OR2_X1 U_g10007B (.ZN(g10007B),.A2(I15210B),.A1(I15209B));
OR2_X1 U_g11267B (.ZN(g11267B),.A2(g11029B),.A1(g11192B));
OR2_X1 U_g11294B (.ZN(g11294B),.A2(g11210B),.A1(g6576B));
OR3_X1 U_g9509B (.ZN(g9509B),.A3(g9111B),.A2(FE_OFN44_g9125B),.A1(g9151B));
OR2_X1 U_g7211B (.ZN(g7211B),.A2(g6067B),.A1(g6647B));
OR2_X1 U_g5404B (.ZN(g5404B),.A2(g3696B),.A1(g4487B));
OR2_X1 U_g4089B (.ZN(g4089B),.A2(I5254B),.A1(g1959B));
OR4_X1 U_I15219B (.ZN(I15219B),.A4(g9833B),.A3(g9936B),.A2(g9907B),.A1(g8172B));
OR2_X1 U_g11219B (.ZN(g11219B),.A2(g11006B),.A1(g11145B));
OR2_X1 U_g6015B (.ZN(g6015B),.A2(g3942B),.A1(g5497B));
OR2_X1 U_g10720B (.ZN(g10720B),.A2(g10667B),.A1(g10304B));
OR2_X1 U_g8265B (.ZN(g8265B),.A2(g4827B),.A1(g7881B));
OR2_X1 U_g5224B (.ZN(g5224B),.A2(g3512B),.A1(g4360B));
OR3_X1 U_g9700B (.ZN(g9700B),.A3(I14827B),.A2(g9667B),.A1(g9358B));
OR2_X1 U_g7106B (.ZN(g7106B),.A2(g5917B),.A1(g6554B));
OR2_X1 U_g8770B (.ZN(g8770B),.A2(g8651B),.A1(g5476B));
OR2_X1 U_g11201B (.ZN(g11201B),.A2(g11011B),.A1(g11152B));
OR3_X1 U_g9950B (.ZN(g9950B),.A3(g9803B),.A2(g9898B),.A1(g9901B));
OR4_X1 U_g9723B (.ZN(g9723B),.A4(I14858B),.A3(g9391B),.A2(g9652B),.A1(g9620B));
OR2_X1 U_g2309B (.ZN(g2309B),.A2(I5358B),.A1(I5357B));
OR2_X1 U_g11266B (.ZN(g11266B),.A2(g11028B),.A1(g11190B));
OR2_X1 U_g10727B (.ZN(g10727B),.A2(g10638B),.A1(g4969B));
OR2_X1 U_g10863B (.ZN(g10863B),.A2(g10750B),.A1(g5531B));
OR2_X1 U_g8429B (.ZN(g8429B),.A2(g8069B),.A1(g8385B));
OR2_X1 U_g9751B (.ZN(g9751B),.A2(g9510B),.A1(g9515B));
OR2_X1 U_g8281B (.ZN(g8281B),.A2(g7818B),.A1(g8097B));
OR2_X1 U_g6910B (.ZN(g6910B),.A2(g5680B),.A1(g6341B));
OR2_X1 U_g8639B (.ZN(g8639B),.A2(g8462B),.A1(g8118B));
OR3_X1 U_g9673B (.ZN(g9673B),.A3(g9274B),.A2(FE_OFN72_g9292B),.A1(g9454B));
OR2_X1 U_g11285B (.ZN(g11285B),.A2(g11161B),.A1(g11255B));
OR2_X1 U_g11305B (.ZN(g11305B),.A2(g11093B),.A1(g11215B));
OR4_X1 U_I15177B (.ZN(I15177B),.A4(g9876B),.A3(g9863B),.A2(g9960B),.A1(g9844B));
OR3_X1 U_g9734B (.ZN(g9734B),.A3(g9426B),.A2(g9428B),.A1(g9415B));
OR3_X1 U_I14827B (.ZN(I14827B),.A3(g9584B),.A2(g9614B),.A1(g9603B));
OR2_X1 U_g5824B (.ZN(g5824B),.A2(g4839B),.A1(g5602B));
OR2_X1 U_g8715B (.ZN(g8715B),.A2(g8687B),.A1(g8416B));
OR2_X1 U_g5762B (.ZN(g5762B),.A2(g5186B),.A1(g5178B));
OR2_X1 U_g6538B (.ZN(g6538B),.A2(g5006B),.A1(g5782B));
OR2_X1 U_g5590B (.ZN(g5590B),.A2(g4723B),.A1(g4718B));
OR2_X1 U_g10726B (.ZN(g10726B),.A2(g10673B),.A1(g10316B));
OR2_X1 U_g3120B (.ZN(g3120B),.A2(I6351B),.A1(I6350B));
OR3_X2 U_g4640B (.ZN(g4640B),.A3(g1527B),.A2(g3563B),.A1(g3348B));
OR2_X1 U_g6093B (.ZN(g6093B),.A2(g4534B),.A1(g5264B));
OR2_X1 U_g8162B (.ZN(g8162B),.A2(g6889B),.A1(g7898B));
OR2_X1 U_g8268B (.ZN(g8268B),.A2(g7613B),.A1(g7962B));
OR2_X1 U_g9569B (.ZN(g9569B),.A2(FE_OFN49_g9030B),.A1(FE_OFN54_g9052B));
OR2_X1 U_g11485B (.ZN(g11485B),.A2(g11462B),.A1(g6646B));
OR2_X1 U_g10797B (.ZN(g10797B),.A2(g10766B),.A1(g6206B));
OR3_X1 U_I14779B (.ZN(I14779B),.A3(g9192B),.A2(g9205B),.A1(g8995B));
OR2_X1 U_g10408B (.ZN(g10408B),.A2(g9097B),.A1(g10298B));
OR2_X1 U_g10635B (.ZN(g10635B),.A2(g7732B),.A1(g10622B));
OR2_X1 U_g2305B (.ZN(g2305B),.A2(I5352B),.A1(I5351B));
OR4_X1 U_I15176B (.ZN(I15176B),.A4(g9836B),.A3(g9897B),.A2(g9908B),.A1(g8176B));
OR2_X1 U_g3435B (.ZN(g3435B),.A2(g2950B),.A1(g2945B));
OR2_X1 U_g9924B (.ZN(g9924B),.A2(g9709B),.A1(g9866B));
OR2_X1 U_g10711B (.ZN(g10711B),.A2(g10690B),.A1(g5547B));
OR2_X1 U_g5814B (.ZN(g5814B),.A2(g4827B),.A1(g5591B));
OR2_X1 U_g5038B (.ZN(g5038B),.A2(g4884B),.A1(g4878B));
OR4_X1 U_I15215B (.ZN(I15215B),.A4(g9879B),.A3(g9854B),.A2(g9965B),.A1(g9840B));
OR2_X1 U_g8226B (.ZN(g8226B),.A2(g7681B),.A1(g7504B));
OR2_X1 U_g7367B (.ZN(g7367B),.A2(g6744B),.A1(g7224B));
OR2_X1 U_g7457B (.ZN(g7457B),.A2(g6404B),.A1(g6873B));
OR2_X1 U_g5229B (.ZN(g5229B),.A2(g3516B),.A1(g4364B));
OR2_X1 U_g5993B (.ZN(g5993B),.A2(g4400B),.A1(g5090B));
OR2_X1 U_g8283B (.ZN(g8283B),.A2(g7820B),.A1(g8098B));
OR2_X1 U_g7971B (.ZN(g7971B),.A2(g7549B),.A1(g5110B));
OR2_X1 U_g8602B (.ZN(g8602B),.A2(g8550B),.A1(g8401B));
OR2_X1 U_g8920B (.ZN(g8920B),.A2(FE_OFN329_g8763B),.A1(g8845B));
OR2_X1 U_g10663B (.ZN(g10663B),.A2(g10581B),.A1(g10237B));
OR2_X1 U_g6074B (.ZN(g6074B),.A2(g1B),.A1(g5349B));
OR2_X1 U_g8261B (.ZN(g8261B),.A2(g3383B),.A1(g7876B));
OR2_X1 U_g10862B (.ZN(g10862B),.A2(g10746B),.A1(g5524B));
OR2_X1 U_g5837B (.ZN(g5837B),.A2(g4224B),.A1(g5640B));
OR2_X1 U_g11333B (.ZN(g11333B),.A2(g11173B),.A1(g11274B));
OR2_X1 U_g6080B (.ZN(g6080B),.A2(g4512B),.A1(g5249B));
OR2_X1 U_g6480B (.ZN(g6480B),.A2(g4971B),.A1(g5721B));
OR2_X1 U_g7740B (.ZN(g7740B),.A2(g6741B),.A1(g7209B));
OR2_X2 U_g10702B (.ZN(g10702B),.A2(g2984B),.A1(g10562B));
OR3_X1 U_g9697B (.ZN(g9697B),.A3(I14822B),.A2(g9606B),.A1(g9665B));
OR2_X1 U_g8203B (.ZN(g8203B),.A2(g7696B),.A1(g7453B));
OR2_X1 U_g9914B (.ZN(g9914B),.A2(g9692B),.A1(g9851B));
OR2_X1 U_g10564B (.ZN(g10564B),.A2(g7368B),.A1(g10560B));
OR2_X1 U_g11484B (.ZN(g11484B),.A2(g11461B),.A1(g6639B));
OR2_X1 U_g5842B (.ZN(g5842B),.A2(g3979B),.A1(g5618B));
OR4_X1 U_I15200B (.ZN(I15200B),.A4(g9880B),.A3(g9848B),.A2(g9962B),.A1(g9837B));
OR2_X1 U_g11609B (.ZN(g11609B),.A2(g11559B),.A1(g11588B));
OR2_X1 U_g8940B (.ZN(g8940B),.A2(FE_OFN332_g8748B),.A1(g8793B));
OR2_X1 U_g11312B (.ZN(g11312B),.A2(g11101B),.A1(g11222B));
OR2_X1 U_g11608B (.ZN(g11608B),.A2(g11558B),.A1(g11587B));
OR2_X1 U_g6000B (.ZN(g6000B),.A2(g3912B),.A1(g5480B));
OR2_X1 U_g8428B (.ZN(g8428B),.A2(g8068B),.A1(g8382B));
OR2_X1 U_g8430B (.ZN(g8430B),.A2(g8070B),.A1(g8386B));
OR2_X1 U_g9922B (.ZN(g9922B),.A2(g9705B),.A1(g9864B));
OR2_X1 U_g8247B (.ZN(g8247B),.A2(g7704B),.A1(g8010B));
OR2_X1 U_g3438B (.ZN(g3438B),.A2(g2944B),.A1(g2939B));
OR4_X1 U_I5576B (.ZN(I5576B),.A4(g444B),.A3(g440B),.A2(g435B),.A1(g431B));
OR2_X1 U_g6924B (.ZN(g6924B),.A2(g4261B),.A1(g6362B));
OR2_X1 U_g5405B (.ZN(g5405B),.A2(FE_OFN221_g3440B),.A1(g4476B));
OR2_X1 U_g8638B (.ZN(g8638B),.A2(g8461B),.A1(g8108B));
OR2_X1 U_g8609B (.ZN(g8609B),.A2(g8555B),.A1(g8408B));
OR2_X1 U_g9995B (.ZN(g9995B),.A2(I15200B),.A1(I15199B));
OR2_X1 U_g8883B (.ZN(g8883B),.A2(FE_OFN329_g8763B),.A1(g8838B));
OR4_X1 U_I15214B (.ZN(I15214B),.A4(g9831B),.A3(g9935B),.A2(g9906B),.A1(g8170B));
OR3_X1 U_g2538B (.ZN(g2538B),.A3(I5649B),.A2(g1458B),.A1(g1466B));
OR2_X1 U_g11329B (.ZN(g11329B),.A2(g11169B),.A1(g11302B));
OR2_X1 U_g4255B (.ZN(g4255B),.A2(g4047B),.A1(g4009B));
OR2_X1 U_g11328B (.ZN(g11328B),.A2(g11168B),.A1(g11299B));
OR3_X1 U_g9704B (.ZN(g9704B),.A3(I14835B),.A2(g9605B),.A1(g9385B));
OR4_X1 U_I5352B (.ZN(I5352B),.A4(g1117B),.A3(g1121B),.A2(g1125B),.A1(g1129B));
OR2_X1 U_g8774B (.ZN(g8774B),.A2(g8654B),.A1(g5499B));
OR3_X1 U_g9954B (.ZN(g9954B),.A3(g9803B),.A2(g9940B),.A1(g9946B));
OR2_X1 U_g10405B (.ZN(g10405B),.A2(g9291B),.A1(g10297B));
OR2_X1 U_g9363B (.ZN(g9363B),.A2(g9192B),.A1(g9205B));
OR2_X1 U_g5849B (.ZN(g5849B),.A2(g4144B),.A1(g4949B));
OR4_X1 U_I5599B (.ZN(I5599B),.A4(g501B),.A3(g506B),.A2(g511B),.A1(g516B));
OR2_X1 U_g7204B (.ZN(g7204B),.A2(I9717B),.A1(g6645B));
OR2_X1 U_g7300B (.ZN(g7300B),.A2(g6326B),.A1(g7139B));
OR2_X1 U_g4293B (.ZN(g4293B),.A2(g4068B),.A1(g4064B));
OR2_X1 U_g9912B (.ZN(g9912B),.A2(g9690B),.A1(g9847B));
OR2_X1 U_g6533B (.ZN(g6533B),.A2(g5002B),.A1(g5771B));
OR2_X1 U_g8816B (.ZN(g8816B),.A2(g8731B),.A1(g7951B));
OR2_X1 U_g9929B (.ZN(g9929B),.A2(g9718B),.A1(g9871B));
OR2_X1 U_g5819B (.ZN(g5819B),.A2(g4876B),.A1(g5625B));
OR3_X1 U_I14831B (.ZN(I14831B),.A3(g9586B),.A2(g9622B),.A1(g9613B));
OR2_X1 U_g5852B (.ZN(g5852B),.A2(g3989B),.A1(g5632B));
OR2_X1 U_g8263B (.ZN(g8263B),.A2(g7720B),.A1(g8032B));
OR2_X1 U_g3431B (.ZN(g3431B),.A2(g2957B),.A1(g2951B));
OR2_X1 U_g8631B (.ZN(g8631B),.A2(g7449B),.A1(g8474B));
OR2_X1 U_g6922B (.ZN(g6922B),.A2(g5694B),.A1(g6352B));
OR2_X1 U_g8817B (.ZN(g8817B),.A2(g8732B),.A1(g7954B));
OR4_X1 U_g9735B (.ZN(g9735B),.A4(g9387B),.A3(g9384B),.A2(g9651B),.A1(g9649B));
OR2_X1 U_g8605B (.ZN(g8605B),.A2(g8553B),.A1(g8404B));
OR2_X1 U_g11263B (.ZN(g11263B),.A2(g11025B),.A1(g11187B));
OR2_X1 U_g6739B (.ZN(g6739B),.A2(g5780B),.A1(g5769B));
OR2_X1 U_g11332B (.ZN(g11332B),.A2(g11172B),.A1(g11273B));
OR2_X1 U_g7143B (.ZN(g7143B),.A2(I9717B),.A1(g6619B));
OR2_X1 U_g6479B (.ZN(g6479B),.A2(g4968B),.A1(g5707B));
OR4_X1 U_I15048B (.ZN(I15048B),.A4(FE_OFN35_g9785B),.A3(FE_OFN61_g9624B),.A2(g9680B),.A1(FE_OFN90_I11360B));
OR2_X1 U_g6501B (.ZN(g6501B),.A2(g4987B),.A1(g5726B));
OR3_X1 U_g9702B (.ZN(g9702B),.A3(I14831B),.A2(g9647B),.A1(g9365B));
OR2_X1 U_g11221B (.ZN(g11221B),.A2(g11007B),.A1(g11146B));
OR3_X1 U_g9952B (.ZN(g9952B),.A3(g9815B),.A2(g9938B),.A1(g9944B));
OR2_X1 U_g11613B (.ZN(g11613B),.A2(g11591B),.A1(g11600B));
OR2_X1 U_g7621B (.ZN(g7621B),.A2(g6994B),.A1(g5108B));
OR2_X1 U_g3399B (.ZN(g3399B),.A2(g2940B),.A1(g2918B));
OR2_X1 U_g11605B (.ZN(g11605B),.A2(g11555B),.A1(g11584B));
OR2_X1 U_g4274B (.ZN(g4274B),.A2(g4058B),.A1(g4054B));
OR3_X1 U_I14602B (.ZN(I14602B),.A3(g9192B),.A2(FE_OFN42_g9205B),.A1(g8995B));
OR4_X1 U_I15033B (.ZN(I15033B),.A4(FE_OFN35_g9785B),.A3(FE_OFN61_g9624B),.A2(FE_OFN33_g9454B),.A1(FE_OFN90_I11360B));
OR2_X1 U_g10717B (.ZN(g10717B),.A2(g10705B),.A1(g6235B));
OR3_X1 U_I5629B (.ZN(I5629B),.A3(g837B),.A2(g841B),.A1(g845B));
OR2_X1 U_g9925B (.ZN(g9925B),.A2(g9712B),.A1(g9867B));
OR2_X1 U_g3819B (.ZN(g3819B),.A2(g9B),.A1(g3275B));
OR2_X1 U_g6912B (.ZN(g6912B),.A2(g4235B),.A1(g6350B));
OR2_X1 U_g10723B (.ZN(g10723B),.A2(g10633B),.A1(g4952B));
OR2_X1 U_g6929B (.ZN(g6929B),.A2(g5704B),.A1(g6360B));
OR2_X1 U_g10646B (.ZN(g10646B),.A2(g7739B),.A1(g10625B));
OR2_X1 U_g9516B (.ZN(g9516B),.A2(FE_OFN44_g9125B),.A1(FE_OFN47_g9151B));
OR2_X1 U_g6626B (.ZN(g6626B),.A2(g123B),.A1(g5934B));
OR4_X1 U_I6350B (.ZN(I6350B),.A4(g2419B),.A3(g2433B),.A2(g2437B),.A1(g2445B));
OR2_X1 U_g11325B (.ZN(g11325B),.A2(g11165B),.A1(g11295B));
OR4_X1 U_I5366B (.ZN(I5366B),.A4(g1296B),.A3(g1292B),.A2(g1284B),.A1(g1280B));
OR3_X1 U_I5649B (.ZN(I5649B),.A3(g1482B),.A2(g1486B),.A1(g1499B));
OR2_X1 U_g6894B (.ZN(g6894B),.A2(g4868B),.A1(g6763B));
OR3_X1 U_g9738B (.ZN(g9738B),.A3(g9506B),.A2(g9447B),.A1(g9417B));
OR2_X1 U_g8383B (.ZN(g8383B),.A2(g5051B),.A1(g8163B));
OR2_X1 U_g8779B (.ZN(g8779B),.A2(g8663B),.A1(g5530B));
OR2_X1 U_g8161B (.ZN(g8161B),.A2(g7185B),.A1(g8005B));
OR2_X2 U_g8451B (.ZN(g8451B),.A2(g8366B),.A1(FE_OFN221_g3440B));
OR2_X1 U_g9915B (.ZN(g9915B),.A2(g9693B),.A1(g9853B));
OR4_X1 U_g2316B (.ZN(g2316B),.A4(I5366B),.A3(g1270B),.A2(g1304B),.A1(g1300B));
OR2_X1 U_g5576B (.ZN(g5576B),.A2(FE_OFN204_g3664B),.A1(g4675B));
OR2_X1 U_g10857B (.ZN(g10857B),.A2(g10738B),.A1(g6090B));
OR2_X1 U_g10793B (.ZN(g10793B),.A2(g10763B),.A1(g6194B));
OR2_X1 U_g7511B (.ZN(g7511B),.A2(g6438B),.A1(g6890B));
OR2_X1 U_g8944B (.ZN(g8944B),.A2(FE_OFN332_g8748B),.A1(g8799B));
OR2_X1 U_g10765B (.ZN(g10765B),.A2(g10680B),.A1(g5492B));
OR2_X1 U_g10549B (.ZN(g10549B),.A2(g10451B),.A1(g4271B));
OR2_X1 U_g7092B (.ZN(g7092B),.A2(g5902B),.A1(g6540B));
OR2_X1 U_g11604B (.ZN(g11604B),.A2(g11554B),.A1(g11583B));
OR2_X1 U_g8434B (.ZN(g8434B),.A2(g8074B),.A1(g8400B));
OR2_X1 U_g6546B (.ZN(g6546B),.A2(g5026B),.A1(g5796B));
OR2_X1 U_g3354B (.ZN(g3354B),.A2(g1216B),.A1(g3121B));
OR2_X1 U_g9928B (.ZN(g9928B),.A2(g9717B),.A1(g9870B));
OR2_X1 U_g11262B (.ZN(g11262B),.A2(g11024B),.A1(g11240B));
OR4_X1 U_g9785B (.ZN(g9785B),.A4(g9363B),.A3(g9388B),.A2(g8995B),.A1(g9010B));
OR2_X1 U_g5867B (.ZN(g5867B),.A2(g4921B),.A1(FE_OFN221_g3440B));
OR2_X1 U_g8210B (.ZN(g8210B),.A2(g7692B),.A1(g7466B));
OR2_X1 U_g10533B (.ZN(g10533B),.A2(g10449B),.A1(g4437B));
OR2_X1 U_g9563B (.ZN(g9563B),.A2(g9030B),.A1(FE_OFN56_g9052B));
OR2_X1 U_g6906B (.ZN(g6906B),.A2(g5674B),.A1(g6791B));
OR2_X1 U_g7375B (.ZN(g7375B),.A2(g6745B),.A1(g7230B));
OR2_X1 U_g7651B (.ZN(g7651B),.A2(FE_OFN350_g3121B),.A1(g7135B));
OR4_X1 U_I5570B (.ZN(I5570B),.A4(g401B),.A3(g406B),.A2(g411B),.A1(g416B));
OR3_X1 U_g9731B (.ZN(g9731B),.A3(g9387B),.A2(g9364B),.A1(g9641B));
OR2_X1 U_g11247B (.ZN(g11247B),.A2(g10949B),.A1(g11097B));
OR4_X1 U_I15045B (.ZN(I15045B),.A4(FE_OFN35_g9785B),.A3(FE_OFN61_g9624B),.A2(g9676B),.A1(FE_OFN90_I11360B));
OR2_X1 U_g10856B (.ZN(g10856B),.A2(g10737B),.A1(g6083B));
OR2_X1 U_g7184B (.ZN(g7184B),.A2(g6047B),.A1(g6625B));
OR2_X1 U_g11612B (.ZN(g11612B),.A2(g11590B),.A1(g11599B));
OR2_X1 U_g7384B (.ZN(g7384B),.A2(g6618B),.A1(g7088B));
OR2_X1 U_g11324B (.ZN(g11324B),.A2(g11164B),.A1(g11271B));
OR2_X1 U_g8922B (.ZN(g8922B),.A2(FE_OFN329_g8763B),.A1(g8822B));
OR4_X1 U_I5358B (.ZN(I5358B),.A4(g1275B),.A3(g1235B),.A2(g1240B),.A1(g1245B));
OR3_X1 U_g9955B (.ZN(g9955B),.A3(g9803B),.A2(g9941B),.A1(g9947B));
OR4_X1 U_g2501B (.ZN(g2501B),.A4(I5576B),.A3(g421B),.A2(g452B),.A1(g448B));
OR2_X1 U_g7231B (.ZN(g7231B),.A2(g6087B),.A1(g6673B));
OR2_X1 U_g6078B (.ZN(g6078B),.A2(g5256B),.A1(g4503B));
OR2_X1 U_g6478B (.ZN(g6478B),.A2(g4967B),.A1(g5706B));
OR2_X1 U_g6907B (.ZN(g6907B),.A2(g5675B),.A1(g6792B));
OR2_X1 U_g6035B (.ZN(g6035B),.A2(g3974B),.A1(g5518B));
OR2_X1 U_g8937B (.ZN(g8937B),.A2(FE_OFN332_g8748B),.A1(g8786B));
OR2_X1 U_g7742B (.ZN(g7742B),.A2(g6743B),.A1(g7217B));
OR2_X1 U_g10722B (.ZN(g10722B),.A2(g10671B),.A1(g10308B));
OR2_X1 U_g9918B (.ZN(g9918B),.A2(g9698B),.A1(g9858B));
OR2_X1 U_g5403B (.ZN(g5403B),.A2(g3695B),.A1(g4486B));
OR2_X1 U_g7926B (.ZN(g7926B),.A2(g6892B),.A1(g7435B));
OR2_X1 U_g6915B (.ZN(g6915B),.A2(g5686B),.A1(g6347B));
OR2_X1 U_g5841B (.ZN(g5841B),.A2(g4230B),.A1(g4914B));
OR4_X1 U_I15220B (.ZN(I15220B),.A4(g9877B),.A3(g9857B),.A2(g9966B),.A1(g9841B));
OR2_X1 U_g10529B (.ZN(g10529B),.A2(I16161B),.A1(I16160B));
OR2_X1 U_g11246B (.ZN(g11246B),.A2(g10948B),.A1(g11094B));
OR2_X1 U_g6002B (.ZN(g6002B),.A2(g4827B),.A1(g5489B));
OR2_X1 U_g7712B (.ZN(g7712B),.A2(FE_OFN350_g3121B),.A1(g7125B));
OR2_X1 U_g8810B (.ZN(g8810B),.A2(g8720B),.A1(g7933B));
OR2_X1 U_g9921B (.ZN(g9921B),.A2(g9703B),.A1(g9862B));
OR2_X1 U_g8432B (.ZN(g8432B),.A2(g8072B),.A1(g8389B));
OR4_X1 U_I15172B (.ZN(I15172B),.A4(g9874B),.A3(g9861B),.A2(g9959B),.A1(g9843B));
OR3_X1 U_I14822B (.ZN(I14822B),.A3(g9582B),.A2(g9604B),.A1(g9597B));
OR2_X1 U_g6928B (.ZN(g6928B),.A2(g5703B),.A1(g6359B));
OR2_X1 U_g8157B (.ZN(g8157B),.A2(g7623B),.A1(FE_OFN192_g6488B));
OR2_X1 U_g6930B (.ZN(g6930B),.A2(g4269B),.A1(g6364B));
OR2_X1 U_g7660B (.ZN(g7660B),.A2(g5867B),.A1(g7059B));
OR2_X1 U_g6899B (.ZN(g6899B),.A2(g32B),.A1(g6463B));
OR2_X1 U_g9392B (.ZN(g9392B),.A2(g9324B),.A1(g9328B));
OR2_X1 U_g11318B (.ZN(g11318B),.A2(g11104B),.A1(g11228B));
OR3_X1 U_I16427B (.ZN(I16427B),.A3(g10382B),.A2(g10383B),.A1(g10683B));
OR2_X1 U_g11227B (.ZN(g11227B),.A2(g11010B),.A1(g11151B));
OR2_X1 U_g11058B (.ZN(g11058B),.A2(g5280B),.A1(g10933B));
OR4_X1 U_I5351B (.ZN(I5351B),.A4(g1133B),.A3(g1137B),.A2(g1141B),.A1(g1145B));
OR3_X1 U_g9708B (.ZN(g9708B),.A3(g9646B),.A2(g9389B),.A1(g9653B));
OR2_X1 U_g6071B (.ZN(g6071B),.A2(g4505B),.A1(g5228B));
OR2_X1 U_g9911B (.ZN(g9911B),.A2(g9689B),.A1(g9846B));
OR2_X1 U_g7102B (.ZN(g7102B),.A2(g5915B),.A1(g6550B));
OR2_X1 U_g7302B (.ZN(g7302B),.A2(g6328B),.A1(g7141B));
OR2_X1 U_g6038B (.ZN(g6038B),.A2(g3979B),.A1(g5528B));
OR2_X1 U_g4239B (.ZN(g4239B),.A2(g4008B),.A1(g4000B));
OR2_X1 U_g8646B (.ZN(g8646B),.A2(g8547B),.A1(g8224B));
OR2_X1 U_g9974B (.ZN(g9974B),.A2(I15177B),.A1(I15176B));
OR2_X1 U_g5823B (.ZN(g5823B),.A2(g4882B),.A1(g5631B));
OR2_X1 U_g6918B (.ZN(g6918B),.A2(g4252B),.A1(g6358B));
OR2_X1 U_g7265B (.ZN(g7265B),.A2(g6204B),.A1(g6756B));
OR4_X1 U_I5804B (.ZN(I5804B),.A4(g2104B),.A3(g2106B),.A2(g2109B),.A1(g2111B));
OR2_X1 U_g5851B (.ZN(g5851B),.A2(g4253B),.A1(g4941B));
OR2_X1 U_g11481B (.ZN(g11481B),.A2(g11458B),.A1(g6624B));
OR2_X1 U_g10336B (.ZN(g10336B),.A2(g9097B),.A1(g10230B));
OR2_X1 U_g7296B (.ZN(g7296B),.A2(g6322B),.A1(g7131B));
OR2_X1 U_g4300B (.ZN(g4300B),.A2(g1212B),.A1(g3546B));
OR2_X1 U_g8647B (.ZN(g8647B),.A2(g8470B),.A1(g8130B));
NAND2_X1 U_g8546B (.ZN(g8546B),.A2(g8390B),.A1(g3983B));
NAND2_X1 U_g2516B (.ZN(g2516B),.A2(I5613B),.A1(I5612B));
NAND2_X1 U_g2987B (.ZN(g2987B),.A2(g883B),.A1(g2481B));
NAND2_X1 U_I5593B (.ZN(I5593B),.A2(I5591B),.A1(g1703B));
NAND2_X1 U_g8970B (.ZN(g8970B),.A2(g8839B),.A1(g5548B));
NAND2_X1 U_I10519B (.ZN(I10519B),.A2(g822B),.A1(g6231B));
NAND2_X1 U_I11279B (.ZN(I11279B),.A2(I11278B),.A1(g305B));
NAND4_X1 U_g7990B (.ZN(g7990B),.A4(g7550B),.A3(g7562B),.A2(FE_OFN80_g2175B),.A1(FE_OFN88_g2178B));
NAND2_X1 U_I11278B (.ZN(I11278B),.A2(g6485B),.A1(g305B));
NAND2_X1 U_g3978B (.ZN(g3978B),.A2(g1822B),.A1(g3207B));
NAND2_X1 U_I5264B (.ZN(I5264B),.A2(I5263B),.A1(g456B));
NAND2_X1 U_I8640B (.ZN(I8640B),.A2(g516B),.A1(g4278B));
NAND2_X1 U_I6761B (.ZN(I6761B),.A2(I6760B),.A1(g2943B));
NAND2_X1 U_I17400B (.ZN(I17400B),.A2(g11416B),.A1(g11418B));
NAND2_X1 U_I5450B (.ZN(I5450B),.A2(I5449B),.A1(g1235B));
NAND2_X1 U_I16060B (.ZN(I16060B),.A2(I16058B),.A1(g10441B));
NAND2_X1 U_I6746B (.ZN(I6746B),.A2(g1453B),.A1(g2938B));
NAND2_X1 U_I11975B (.ZN(I11975B),.A2(I11973B),.A1(g1462B));
NAND2_X1 U_I12136B (.ZN(I12136B),.A2(g131B),.A1(g6038B));
NAND2_X1 U_I11937B (.ZN(I11937B),.A2(I11935B),.A1(g1458B));
NAND2_X1 U_g2959B (.ZN(g2959B),.A2(I6168B),.A1(I6167B));
NAND2_X1 U_I5878B (.ZN(I5878B),.A2(g2115B),.A1(g2120B));
NAND2_X1 U_g2517B (.ZN(g2517B),.A2(I5620B),.A1(I5619B));
NAND2_X1 U_g5552B (.ZN(g5552B),.A2(FE_OFN223_g4401B),.A1(g4777B));
NAND2_X1 U_I6468B (.ZN(I6468B),.A2(I6467B),.A1(g23B));
NAND2_X1 U_I8796B (.ZN(I8796B),.A2(I8795B),.A1(g4672B));
NAND2_X1 U_g10392B (.ZN(g10392B),.A2(I15892B),.A1(I15891B));
NAND2_X1 U_I5611B (.ZN(I5611B),.A2(g1284B),.A1(g1280B));
NAND2_X1 U_g8738B (.ZN(g8738B),.A2(FE_OFN200_g4921B),.A1(g8688B));
NAND2_X1 U_I6716B (.ZN(I6716B),.A2(I6714B),.A1(g201B));
NAND2_X1 U_g2310B (.ZN(g2310B),.A2(g605B),.A1(g591B));
NAND2_X1 U_I7685B (.ZN(I7685B),.A2(I7683B),.A1(g3460B));
NAND2_X1 U_g3056B (.ZN(g3056B),.A2(g599B),.A1(g2374B));
NAND2_X1 U_I12108B (.ZN(I12108B),.A2(I12106B),.A1(g135B));
NAND3_X1 U_g3529B (.ZN(g3529B),.A3(g2325B),.A2(g3062B),.A1(g2310B));
NAND2_X1 U_I6747B (.ZN(I6747B),.A2(I6746B),.A1(g2938B));
NAND2_X1 U_g2236B (.ZN(g2236B),.A2(I5231B),.A1(I5230B));
NAND2_X1 U_g7584B (.ZN(g7584B),.A2(I12076B),.A1(I12075B));
NAND2_X1 U_I15870B (.ZN(I15870B),.A2(FE_OFN239_g1796B),.A1(g10291B));
NAND2_X1 U_I16067B (.ZN(I16067B),.A2(I16065B),.A1(FE_OFN237_g1806B));
NAND2_X1 U_I7562B (.ZN(I7562B),.A2(g654B),.A1(g3533B));
NAND2_X1 U_I13531B (.ZN(I13531B),.A2(I13529B),.A1(g8253B));
NAND2_X1 U_I8797B (.ZN(I8797B),.A2(I8795B),.A1(g1145B));
NAND2_X1 U_I17584B (.ZN(I17584B),.A2(g11515B),.A1(g11217B));
NAND2_X1 U_I11936B (.ZN(I11936B),.A2(I11935B),.A1(g5857B));
NAND2_X1 U_I15257B (.ZN(I15257B),.A2(I15256B),.A1(g9974B));
NAND2_X1 U_g8402B (.ZN(g8402B),.A2(I13506B),.A1(I13505B));
NAND3_X1 U_g8824B (.ZN(g8824B),.A3(g8512B),.A2(g8501B),.A1(g8502B));
NAND2_X1 U_I6186B (.ZN(I6186B),.A2(g466B),.A1(g2511B));
NAND2_X1 U_g11496B (.ZN(g11496B),.A2(I17505B),.A1(I17504B));
NAND2_X1 U_I16001B (.ZN(I16001B),.A2(I15999B),.A1(FE_OFN247_g1771B));
NAND2_X1 U_I6125B (.ZN(I6125B),.A2(I6124B),.A1(g2215B));
NAND2_X1 U_I11909B (.ZN(I11909B),.A2(I11907B),.A1(g1474B));
NAND2_X1 U_I12040B (.ZN(I12040B),.A2(I12038B),.A1(g1466B));
NAND2_X1 U_I13909B (.ZN(I13909B),.A2(I13907B),.A1(g1432B));
NAND2_X1 U_g3625B (.ZN(g3625B),.A2(I6772B),.A1(I6771B));
NAND2_X1 U_I11908B (.ZN(I11908B),.A2(I11907B),.A1(g5838B));
NAND2_X1 U_g10470B (.ZN(g10470B),.A2(I16009B),.A1(I16008B));
NAND2_X1 U_I13908B (.ZN(I13908B),.A2(I13907B),.A1(g8265B));
NAND2_X1 U_g3813B (.ZN(g3813B),.A2(I7035B),.A1(I7034B));
NAND2_X1 U_I8650B (.ZN(I8650B),.A2(g778B),.A1(g4824B));
NAND2_X1 U_g6207B (.ZN(g6207B),.A2(I9948B),.A1(I9947B));
NAND2_X1 U_I16066B (.ZN(I16066B),.A2(I16065B),.A1(g10428B));
NAND2_X1 U_g2948B (.ZN(g2948B),.A2(I6145B),.A1(I6144B));
NAND2_X1 U_I11242B (.ZN(I11242B),.A2(I11241B),.A1(g6760B));
NAND2_X1 U_g10467B (.ZN(g10467B),.A2(I15994B),.A1(I15993B));
NAND2_X1 U_I6187B (.ZN(I6187B),.A2(I6186B),.A1(g2511B));
NAND2_X1 U_g6488B (.ZN(g6488B),.A2(g6019B),.A1(g6027B));
NAND2_X1 U_I5500B (.ZN(I5500B),.A2(g1007B),.A1(g1255B));
NAND2_X1 U_I11974B (.ZN(I11974B),.A2(I11973B),.A1(g5852B));
NAND2_X1 U_I12062B (.ZN(I12062B),.A2(I12060B),.A1(g1478B));
NAND2_X1 U_g5300B (.ZN(g5300B),.A2(I8772B),.A1(I8771B));
NAND2_X1 U_I5184B (.ZN(I5184B),.A2(g1515B),.A1(g1415B));
NAND2_X1 U_I13293B (.ZN(I13293B),.A2(g8161B),.A1(g1882B));
NAND2_X1 U_I6200B (.ZN(I6200B),.A2(I6199B),.A1(g2525B));
NAND2_X1 U_I13265B (.ZN(I13265B),.A2(g8154B),.A1(g1909B));
NAND2_X1 U_I5024B (.ZN(I5024B),.A2(I5023B),.A1(g995B));
NAND2_X1 U_I7863B (.ZN(I7863B),.A2(g774B),.A1(g4099B));
NAND2_X1 U_g8705B (.ZN(g8705B),.A2(I13992B),.A1(I13991B));
NAND2_X1 U_g8471B (.ZN(g8471B),.A2(I13661B),.A1(I13660B));
NAND2_X1 U_I15256B (.ZN(I15256B),.A2(g9968B),.A1(g9974B));
NAND2_X1 U_I6145B (.ZN(I6145B),.A2(I6143B),.A1(g646B));
NAND2_X1 U_I13992B (.ZN(I13992B),.A2(I13990B),.A1(g8688B));
NAND2_X1 U_I11510B (.ZN(I11510B),.A2(I11508B),.A1(FE_OFN237_g1806B));
NAND2_X1 U_g10853B (.ZN(g10853B),.A2(g5034B),.A1(g10731B));
NAND2_X1 U_I5231B (.ZN(I5231B),.A2(I5229B),.A1(g148B));
NAND2_X1 U_I12047B (.ZN(I12047B),.A2(I12045B),.A1(g1486B));
NAND2_X1 U_I10771B (.ZN(I10771B),.A2(I10769B),.A1(g1801B));
NAND2_X1 U_g10477B (.ZN(g10477B),.A2(I16046B),.A1(I16045B));
NAND2_X1 U_g7582B (.ZN(g7582B),.A2(I12062B),.A1(I12061B));
NAND2_X1 U_I5104B (.ZN(I5104B),.A2(g435B),.A1(g431B));
NAND2_X1 U_g8409B (.ZN(g8409B),.A2(I13531B),.A1(I13530B));
NAND2_X1 U_I6447B (.ZN(I6447B),.A2(FE_OFN236_g1776B),.A1(g2264B));
NAND2_X1 U_I4956B (.ZN(I4956B),.A2(I4954B),.A1(g327B));
NAND2_X1 U_I5613B (.ZN(I5613B),.A2(I5611B),.A1(g1284B));
NAND2_X1 U_I8481B (.ZN(I8481B),.A2(I8479B),.A1(g3530B));
NAND2_X1 U_g5278B (.ZN(g5278B),.A2(I8740B),.A1(I8739B));
NAND2_X1 U_I6880B (.ZN(I6880B),.A2(I6879B),.A1(g3301B));
NAND2_X1 U_I15431B (.ZN(I15431B),.A2(I15430B),.A1(g10001B));
NAND2_X1 U_g5548B (.ZN(g5548B),.A2(FE_OFN223_g4401B),.A1(g1840B));
NAND4_X1 U_g7671B (.ZN(g7671B),.A4(FE_OFN96_g2169B),.A3(FE_OFN91_g2172B),.A2(g2175B),.A1(g2178B));
NAND2_X1 U_I12020B (.ZN(I12020B),.A2(I12019B),.A1(g6049B));
NAND2_X1 U_g10665B (.ZN(g10665B),.A2(I16332B),.A1(I16331B));
NAND2_X1 U_I16469B (.ZN(I16469B),.A2(I16467B),.A1(g10518B));
NAND2_X1 U_I5014B (.ZN(I5014B),.A2(I5013B),.A1(g1007B));
NAND2_X1 U_I13523B (.ZN(I13523B),.A2(I13521B),.A1(g8249B));
NAND2_X1 U_I16039B (.ZN(I16039B),.A2(I16037B),.A1(FE_OFN252_g1791B));
NAND2_X1 U_I16468B (.ZN(I16468B),.A2(I16467B),.A1(g10716B));
NAND2_X1 U_I12046B (.ZN(I12046B),.A2(I12045B),.A1(g5814B));
NAND2_X1 U_g4476B (.ZN(g4476B),.A2(g3071B),.A1(g3807B));
NAND2_X1 U_g10476B (.ZN(g10476B),.A2(I16039B),.A1(I16038B));
NAND2_X1 U_I16038B (.ZN(I16038B),.A2(I16037B),.A1(g10363B));
NAND2_X1 U_I8676B (.ZN(I8676B),.A2(g1027B),.A1(g4374B));
NAND2_X1 U_I12113B (.ZN(I12113B),.A2(g162B),.A1(g6002B));
NAND2_X1 U_I8761B (.ZN(I8761B),.A2(g1129B),.A1(g4616B));
NAND2_X1 U_g3204B (.ZN(g3204B),.A2(g2061B),.A1(g2571B));
NAND2_X1 U_I15993B (.ZN(I15993B),.A2(I15992B),.A1(g10430B));
NAND2_X1 U_I5036B (.ZN(I5036B),.A2(I5034B),.A1(g1019B));
NAND2_X1 U_I14263B (.ZN(I14263B),.A2(g1814B),.A1(g8843B));
NAND2_X1 U_g8298B (.ZN(g8298B),.A2(I13250B),.A1(I13249B));
NAND2_X1 U_I5135B (.ZN(I5135B),.A2(g525B),.A1(g521B));
NAND2_X1 U_g2405B (.ZN(g2405B),.A2(I5486B),.A1(I5485B));
NAND2_X1 U_I7034B (.ZN(I7034B),.A2(I7033B),.A1(g3089B));
NAND2_X1 U_I15443B (.ZN(I15443B),.A2(I15441B),.A1(g10007B));
NAND2_X1 U_I6166B (.ZN(I6166B),.A2(g153B),.A1(g2236B));
NAND2_X1 U_I8624B (.ZN(I8624B),.A2(g511B),.A1(g4267B));
NAND2_X1 U_I16015B (.ZN(I16015B),.A2(g1781B),.A1(g10441B));
NAND2_X1 U_I8677B (.ZN(I8677B),.A2(I8676B),.A1(g4374B));
NAND2_X1 U_I8576B (.ZN(I8576B),.A2(I8575B),.A1(g4234B));
NAND2_X1 U_I14613B (.ZN(I14613B),.A2(I14612B),.A1(g9204B));
NAND2_X1 U_I8716B (.ZN(I8716B),.A2(I8715B),.A1(g4601B));
NAND2_X1 U_g3530B (.ZN(g3530B),.A2(I6716B),.A1(I6715B));
NAND2_X1 U_g8405B (.ZN(g8405B),.A2(I13515B),.A1(I13514B));
NAND4_X1 U_g4104B (.ZN(g4104B),.A4(g3200B),.A3(g2439B),.A2(g3247B),.A1(g3215B));
NAND2_X1 U_I12003B (.ZN(I12003B),.A2(I12002B),.A1(g5996B));
NAND2_X1 U_g2177B (.ZN(g2177B),.A2(I5128B),.A1(I5127B));
NAND2_X1 U_g3010B (.ZN(g3010B),.A2(g2399B),.A1(g2382B));
NAND2_X1 U_g5179B (.ZN(g5179B),.A2(I8577B),.A1(I8576B));
NAND2_X1 U_I17395B (.ZN(I17395B),.A2(I17393B),.A1(g11414B));
NAND2_X1 U_g7067B (.ZN(g7067B),.A2(I11280B),.A1(I11279B));
NAND4_X1 U_g7994B (.ZN(g7994B),.A4(g7550B),.A3(FE_OFN91_g2172B),.A2(g7574B),.A1(FE_OFN88_g2178B));
NAND2_X1 U_I6167B (.ZN(I6167B),.A2(I6166B),.A1(g2236B));
NAND2_X1 U_I5265B (.ZN(I5265B),.A2(I5263B),.A1(g461B));
NAND2_X1 U_I6989B (.ZN(I6989B),.A2(I6988B),.A1(g2760B));
NAND2_X1 U_I13274B (.ZN(I13274B),.A2(I13272B),.A1(g8158B));
NAND2_X1 U_I10507B (.ZN(I10507B),.A2(g786B),.A1(g6221B));
NAND2_X1 U_I13530B (.ZN(I13530B),.A2(I13529B),.A1(g704B));
NAND2_X1 U_I5164B (.ZN(I5164B),.A2(g1499B),.A1(g1508B));
NAND2_X1 U_g9107B (.ZN(g9107B),.A2(I14444B),.A1(I14443B));
NAND2_X1 U_I9559B (.ZN(I9559B),.A2(I9557B),.A1(g782B));
NAND2_X1 U_I8577B (.ZN(I8577B),.A2(I8575B),.A1(g496B));
NAND2_X1 U_g2510B (.ZN(g2510B),.A2(I5593B),.A1(I5592B));
NAND2_X1 U_g8177B (.ZN(g8177B),.A2(I13078B),.A1(I13077B));
NAND2_X1 U_I8717B (.ZN(I8717B),.A2(I8715B),.A1(g4052B));
NAND2_X1 U_I5296B (.ZN(I5296B),.A2(I5295B),.A1(g794B));
NAND2_X1 U_g5209B (.ZN(g5209B),.A2(I8626B),.A1(I8625B));
NAND4_X1 U_g7950B (.ZN(g7950B),.A4(FE_OFN96_g2169B),.A3(g7562B),.A2(g7574B),.A1(g6941B));
NAND2_X1 U_g2088B (.ZN(g2088B),.A2(I4912B),.A1(I4911B));
NAND2_X1 U_I16000B (.ZN(I16000B),.A2(I15999B),.A1(g10432B));
NAND2_X1 U_I5371B (.ZN(I5371B),.A2(g976B),.A1(g971B));
NAND2_X1 U_g2215B (.ZN(g2215B),.A2(I5186B),.A1(I5185B));
NAND2_X1 U_g7101B (.ZN(g7101B),.A2(g2364B),.A1(g6617B));
NAND2_X1 U_I5675B (.ZN(I5675B),.A2(g1223B),.A1(g1218B));
NAND2_X1 U_I8544B (.ZN(I8544B),.A2(I8543B),.A1(g4218B));
NAND2_X1 U_g6577B (.ZN(g6577B),.A2(I10521B),.A1(I10520B));
NAND2_X1 U_I5297B (.ZN(I5297B),.A2(I5295B),.A1(g798B));
NAND2_X1 U_I13537B (.ZN(I13537B),.A2(g8157B),.A1(g658B));
NAND2_X1 U_I13283B (.ZN(I13283B),.A2(g8159B),.A1(g1927B));
NAND2_X1 U_g4749B (.ZN(g4749B),.A2(g2061B),.A1(g3710B));
NAND2_X1 U_I11982B (.ZN(I11982B),.A2(I11980B),.A1(g1482B));
NAND2_X1 U_I8514B (.ZN(I8514B),.A2(I8513B),.A1(g4873B));
NAND2_X1 U_I13091B (.ZN(I13091B),.A2(I13089B),.A1(g1840B));
NAND2_X1 U_g2943B (.ZN(g2943B),.A2(I6126B),.A1(I6125B));
NAND2_X1 U_I15908B (.ZN(I15908B),.A2(I15906B),.A1(g10302B));
NAND2_X1 U_I6879B (.ZN(I6879B),.A2(g1351B),.A1(g3301B));
NAND2_X1 U_I8763B (.ZN(I8763B),.A2(I8761B),.A1(g1129B));
NAND2_X1 U_I5449B (.ZN(I5449B),.A2(g991B),.A1(g1235B));
NAND3_X1 U_g8825B (.ZN(g8825B),.A3(g8506B),.A2(g8738B),.A1(g8502B));
NAND2_X1 U_I16007B (.ZN(I16007B),.A2(FE_OFN236_g1776B),.A1(g10434B));
NAND2_X1 U_I5865B (.ZN(I5865B),.A2(g2105B),.A1(g2107B));
NAND2_X1 U_I5604B (.ZN(I5604B),.A2(g1153B),.A1(g1149B));
NAND2_X1 U_g2433B (.ZN(g2433B),.A2(I5518B),.A1(I5517B));
NAND2_X1 U_I6111B (.ZN(I6111B),.A2(I6109B),.A1(g1494B));
NAND2_X1 U_g2096B (.ZN(g2096B),.A2(I4930B),.A1(I4929B));
NAND2_X1 U_I13522B (.ZN(I13522B),.A2(I13521B),.A1(g695B));
NAND2_X1 U_I10770B (.ZN(I10770B),.A2(I10769B),.A1(g5944B));
NAND2_X1 U_g6027B (.ZN(g6027B),.A2(FE_OFN200_g4921B),.A1(g4566B));
NAND4_X1 U_g7992B (.ZN(g7992B),.A4(FE_OFN96_g2169B),.A3(FE_OFN91_g2172B),.A2(g7574B),.A1(FE_OFN88_g2178B));
NAND2_X1 U_I5539B (.ZN(I5539B),.A2(I5538B),.A1(g1270B));
NAND2_X1 U_I17394B (.ZN(I17394B),.A2(I17393B),.A1(g11415B));
NAND2_X1 U_I13553B (.ZN(I13553B),.A2(I13552B),.A1(g668B));
NAND2_X1 U_I8642B (.ZN(I8642B),.A2(I8640B),.A1(g516B));
NAND2_X1 U_g7573B (.ZN(g7573B),.A2(I12047B),.A1(I12046B));
NAND2_X1 U_g11416B (.ZN(g11416B),.A2(I17297B),.A1(I17296B));
NAND2_X1 U_g6003B (.ZN(g6003B),.A2(g5548B),.A1(g5552B));
NAND2_X1 U_g8934B (.ZN(g8934B),.A2(I14279B),.A1(I14278B));
NAND2_X1 U_I15992B (.ZN(I15992B),.A2(g2677B),.A1(g10430B));
NAND2_X1 U_I7683B (.ZN(I7683B),.A2(g3460B),.A1(g1023B));
NAND2_X1 U_I4910B (.ZN(I4910B),.A2(g318B),.A1(g386B));
NAND4_X1 U_g3209B (.ZN(g3209B),.A4(g2571B),.A3(g2564B),.A2(g2061B),.A1(g2550B));
NAND2_X1 U_I6794B (.ZN(I6794B),.A2(I6792B),.A1(g143B));
NAND2_X1 U_I10521B (.ZN(I10521B),.A2(I10519B),.A1(g822B));
NAND2_X1 U_I5486B (.ZN(I5486B),.A2(I5484B),.A1(g1011B));
NAND2_X1 U_I15442B (.ZN(I15442B),.A2(I15441B),.A1(g10013B));
NAND2_X1 U_g6858B (.ZN(g6858B),.A2(I10932B),.A1(I10931B));
NAND2_X1 U_I5185B (.ZN(I5185B),.A2(I5184B),.A1(g1415B));
NAND2_X1 U_g5304B (.ZN(g5304B),.A2(I8780B),.A1(I8779B));
NAND2_X1 U_g2354B (.ZN(g2354B),.A2(g1520B),.A1(g1515B));
NAND2_X1 U_I15615B (.ZN(I15615B),.A2(g10153B),.A1(g10043B));
NAND2_X1 U_I17281B (.ZN(I17281B),.A2(g11219B),.A1(g11221B));
NAND2_X1 U_I5470B (.ZN(I5470B),.A2(I5468B),.A1(g999B));
NAND2_X1 U_I11509B (.ZN(I11509B),.A2(I11508B),.A1(g6580B));
NAND2_X1 U_I5025B (.ZN(I5025B),.A2(I5023B),.A1(g1275B));
NAND2_X1 U_I11508B (.ZN(I11508B),.A2(g1806B),.A1(g6580B));
NAND2_X1 U_I15430B (.ZN(I15430B),.A2(g9995B),.A1(g10001B));
NAND2_X1 U_I14612B (.ZN(I14612B),.A2(g611B),.A1(g9204B));
NAND2_X1 U_g4675B (.ZN(g4675B),.A2(g3247B),.A1(g4073B));
NAND2_X1 U_I14272B (.ZN(I14272B),.A2(I14270B),.A1(g1822B));
NAND2_X1 U_g2979B (.ZN(g2979B),.A2(I6209B),.A1(I6208B));
NAND2_X1 U_I17290B (.ZN(I17290B),.A2(I17288B),.A1(g11223B));
NAND2_X1 U_g5269B (.ZN(g5269B),.A2(I8717B),.A1(I8716B));
NAND2_X1 U_g4297B (.ZN(g4297B),.A2(I7564B),.A1(I7563B));
NAND2_X1 U_I12002B (.ZN(I12002B),.A2(g153B),.A1(g5996B));
NAND2_X1 U_I5006B (.ZN(I5006B),.A2(I5005B),.A1(g421B));
NAND2_X1 U_I12128B (.ZN(I12128B),.A2(I12126B),.A1(g170B));
NAND2_X1 U_I5105B (.ZN(I5105B),.A2(I5104B),.A1(g431B));
NAND2_X1 U_I6323B (.ZN(I6323B),.A2(I6322B),.A1(g2050B));
NAND2_X1 U_g7588B (.ZN(g7588B),.A2(I12094B),.A1(I12093B));
NAND2_X1 U_I6666B (.ZN(I6666B),.A2(I6664B),.A1(g2776B));
NAND2_X1 U_g3623B (.ZN(g3623B),.A2(I6762B),.A1(I6761B));
NAND2_X1 U_I5373B (.ZN(I5373B),.A2(I5371B),.A1(g976B));
NAND2_X1 U_I8529B (.ZN(I8529B),.A2(I8527B),.A1(g481B));
NAND2_X1 U_I5283B (.ZN(I5283B),.A2(I5282B),.A1(g758B));
NAND2_X1 U_I7224B (.ZN(I7224B),.A2(I7223B),.A1(g2981B));
NAND2_X1 U_I5007B (.ZN(I5007B),.A2(I5005B),.A1(g312B));
NAND2_X1 U_I5459B (.ZN(I5459B),.A2(g1003B),.A1(g1240B));
NAND2_X1 U_I17297B (.ZN(I17297B),.A2(I17295B),.A1(g11227B));
NAND3_X1 U_g8746B (.ZN(g8746B),.A3(g46B),.A2(g47B),.A1(g8617B));
NAND2_X1 U_I6143B (.ZN(I6143B),.A2(g646B),.A1(g1976B));
NAND2_X1 U_I5015B (.ZN(I5015B),.A2(I5013B),.A1(g1011B));
NAND2_X1 U_g8932B (.ZN(g8932B),.A2(I14265B),.A1(I14264B));
NAND2_X1 U_I16073B (.ZN(I16073B),.A2(I16072B),.A1(g845B));
NAND2_X1 U_I6988B (.ZN(I6988B),.A2(g986B),.A1(g2760B));
NAND2_X1 U_g3205B (.ZN(g3205B),.A2(g2571B),.A1(g1814B));
NAND2_X1 U_I8652B (.ZN(I8652B),.A2(I8650B),.A1(g778B));
NAND2_X1 U_I9558B (.ZN(I9558B),.A2(I9557B),.A1(g5598B));
NAND2_X1 U_I5203B (.ZN(I5203B),.A2(I5202B),.A1(g369B));
NAND2_X1 U_g7533B (.ZN(g7533B),.A2(I11937B),.A1(I11936B));
NAND2_X1 U_g3634B (.ZN(g3634B),.A2(I6807B),.A1(I6806B));
NAND2_X1 U_I6792B (.ZN(I6792B),.A2(g143B),.A1(g2959B));
NAND2_X1 U_g3304B (.ZN(g3304B),.A2(I6469B),.A1(I6468B));
NAND2_X1 U_I12145B (.ZN(I12145B),.A2(I12143B),.A1(g158B));
NAND2_X1 U_g7596B (.ZN(g7596B),.A2(I12128B),.A1(I12127B));
NAND2_X1 U_I13302B (.ZN(I13302B),.A2(I13300B),.A1(g8162B));
NAND2_X1 U_I5502B (.ZN(I5502B),.A2(I5500B),.A1(g1007B));
NAND2_X1 U_I9574B (.ZN(I9574B),.A2(g818B),.A1(g5608B));
NAND2_X1 U_g3273B (.ZN(g3273B),.A2(I6449B),.A1(I6448B));
NAND2_X1 U_I8670B (.ZN(I8670B),.A2(I8669B),.A1(g4831B));
NAND2_X1 U_I7035B (.ZN(I7035B),.A2(I7033B),.A1(g1868B));
NAND2_X1 U_I15453B (.ZN(I15453B),.A2(I15451B),.A1(g10019B));
NAND2_X1 U_I8625B (.ZN(I8625B),.A2(I8624B),.A1(g4267B));
NAND2_X1 U_I7876B (.ZN(I7876B),.A2(I7875B),.A1(g4109B));
NAND2_X1 U_I14203B (.ZN(I14203B),.A2(I14202B),.A1(g8825B));
NAND2_X1 U_I15607B (.ZN(I15607B),.A2(g10144B),.A1(g10149B));
NAND2_X1 U_g2274B (.ZN(g2274B),.A2(I5325B),.A1(I5324B));
NAND2_X1 U_I8740B (.ZN(I8740B),.A2(I8738B),.A1(g1121B));
NAND2_X1 U_I17296B (.ZN(I17296B),.A2(I17295B),.A1(g11229B));
NAND2_X1 U_g10507B (.ZN(g10507B),.A2(g5859B),.A1(g10434B));
NAND2_X1 U_g2325B (.ZN(g2325B),.A2(g617B),.A1(g611B));
NAND2_X1 U_I8606B (.ZN(I8606B),.A2(I8604B),.A1(g506B));
NAND2_X1 U_I12087B (.ZN(I12087B),.A2(I12085B),.A1(g1470B));
NAND2_X1 U_I13249B (.ZN(I13249B),.A2(I13248B),.A1(g1891B));
NAND2_X1 U_I13248B (.ZN(I13248B),.A2(g8148B),.A1(g1891B));
NAND2_X1 U_I13552B (.ZN(I13552B),.A2(g8262B),.A1(g668B));
NAND2_X1 U_g2106B (.ZN(g2106B),.A2(I4980B),.A1(I4979B));
NAND2_X1 U_I12069B (.ZN(I12069B),.A2(I12067B),.A1(g139B));
NAND2_X1 U_g9204B (.ZN(g9204B),.A2(g8942B),.A1(g6019B));
NAND2_X1 U_I12068B (.ZN(I12068B),.A2(I12067B),.A1(g6045B));
NAND2_X1 U_I17503B (.ZN(I17503B),.A2(g5269B),.A1(g11430B));
NAND2_X1 U_I7877B (.ZN(I7877B),.A2(I7875B),.A1(g810B));
NAND2_X1 U_I5165B (.ZN(I5165B),.A2(I5164B),.A1(g1508B));
NAND2_X1 U_g6740B (.ZN(g6740B),.A2(g2550B),.A1(g6131B));
NAND2_X1 U_I6289B (.ZN(I6289B),.A2(I6287B),.A1(g981B));
NAND2_X1 U_I6777B (.ZN(I6777B),.A2(g650B),.A1(g2892B));
NAND2_X1 U_g5171B (.ZN(g5171B),.A2(I8563B),.A1(I8562B));
NAND2_X1 U_I15891B (.ZN(I15891B),.A2(I15890B),.A1(g853B));
NAND2_X1 U_I13090B (.ZN(I13090B),.A2(I13089B),.A1(g8006B));
NAND2_X1 U_g11474B (.ZN(g11474B),.A2(I17461B),.A1(I17460B));
NAND4_X1 U_g7942B (.ZN(g7942B),.A4(g7550B),.A3(g7562B),.A2(FE_OFN80_g2175B),.A1(g6941B));
NAND2_X1 U_I5538B (.ZN(I5538B),.A2(g1023B),.A1(g1270B));
NAND2_X1 U_I7563B (.ZN(I7563B),.A2(I7562B),.A1(g3533B));
NAND2_X1 U_I13513B (.ZN(I13513B),.A2(g8248B),.A1(g686B));
NAND2_X1 U_g2107B (.ZN(g2107B),.A2(I4987B),.A1(I4986B));
NAND2_X1 U_g2223B (.ZN(g2223B),.A2(I5204B),.A1(I5203B));
NAND2_X1 U_I13505B (.ZN(I13505B),.A2(I13504B),.A1(g677B));
NAND2_X1 U_I6209B (.ZN(I6209B),.A2(I6207B),.A1(g802B));
NAND2_X1 U_I12086B (.ZN(I12086B),.A2(I12085B),.A1(g5842B));
NAND2_X1 U_I8545B (.ZN(I8545B),.A2(I8543B),.A1(g486B));
NAND2_X1 U_I8180B (.ZN(I8180B),.A2(I8178B),.A1(FE_OFN253_g1786B));
NAND2_X1 U_g2115B (.ZN(g2115B),.A2(I5015B),.A1(I5014B));
NAND2_X1 U_I8591B (.ZN(I8591B),.A2(I8589B),.A1(g501B));
NAND2_X1 U_I10931B (.ZN(I10931B),.A2(I10930B),.A1(g5863B));
NAND2_X1 U_I17402B (.ZN(I17402B),.A2(I17400B),.A1(g11416B));
NAND2_X1 U_g8307B (.ZN(g8307B),.A2(I13295B),.A1(I13294B));
NAND2_X1 U_I12144B (.ZN(I12144B),.A2(I12143B),.A1(g6000B));
NAND2_X1 U_I10520B (.ZN(I10520B),.A2(I10519B),.A1(g6231B));
NAND2_X1 U_I5263B (.ZN(I5263B),.A2(FE_OFN254_g461B),.A1(g456B));
NAND2_X1 U_g8757B (.ZN(g8757B),.A2(FE_OFN223_g4401B),.A1(g8599B));
NAND2_X1 U_I6714B (.ZN(I6714B),.A2(g201B),.A1(g2961B));
NAND2_X1 U_I14211B (.ZN(I14211B),.A2(I14209B),.A1(g599B));
NAND2_X1 U_I8515B (.ZN(I8515B),.A2(I8513B),.A1(g3513B));
NAND2_X1 U_g2272B (.ZN(g2272B),.A2(I5317B),.A1(I5316B));
NAND2_X1 U_I9946B (.ZN(I9946B),.A2(g1796B),.A1(g5233B));
NAND2_X1 U_I8750B (.ZN(I8750B),.A2(g1125B),.A1(g4613B));
NAND2_X1 U_I5605B (.ZN(I5605B),.A2(I5604B),.A1(g1149B));
NAND2_X1 U_g8880B (.ZN(g8880B),.A2(I14204B),.A1(I14203B));
NAND2_X1 U_I16051B (.ZN(I16051B),.A2(g10434B),.A1(g837B));
NAND2_X1 U_I16072B (.ZN(I16072B),.A2(g10438B),.A1(g845B));
NAND2_X1 U_g10440B (.ZN(g10440B),.A2(g6037B),.A1(g10360B));
NAND2_X1 U_g8612B (.ZN(g8612B),.A2(I13859B),.A1(I13858B));
NAND2_X1 U_I15872B (.ZN(I15872B),.A2(I15870B),.A1(FE_OFN239_g1796B));
NAND2_X1 U_I8528B (.ZN(I8528B),.A2(I8527B),.A1(g4879B));
NAND2_X1 U_g8629B (.ZN(g8629B),.A2(I13902B),.A1(I13901B));
NAND4_X1 U_g8542B (.ZN(g8542B),.A4(g8390B),.A3(g1814B),.A2(g1828B),.A1(g2571B));
NAND2_X1 U_I9947B (.ZN(I9947B),.A2(I9946B),.A1(g5233B));
NAND2_X1 U_I6838B (.ZN(I6838B),.A2(I6836B),.A1(g806B));
NAND2_X1 U_g7583B (.ZN(g7583B),.A2(I12069B),.A1(I12068B));
NAND2_X1 U_g4803B (.ZN(g4803B),.A2(FE_OFN325_g18B),.A1(g3664B));
NAND2_X1 U_I17307B (.ZN(I17307B),.A2(I17305B),.A1(g11231B));
NAND2_X1 U_g4538B (.ZN(g4538B),.A2(g2399B),.A1(g3475B));
NAND2_X1 U_I15452B (.ZN(I15452B),.A2(I15451B),.A1(g10025B));
NAND2_X1 U_I13857B (.ZN(I13857B),.A2(g1448B),.A1(g8270B));
NAND2_X1 U_I14202B (.ZN(I14202B),.A2(g591B),.A1(g8825B));
NAND2_X1 U_I13765B (.ZN(I13765B),.A2(g8417B),.A1(g731B));
NAND2_X1 U_g2260B (.ZN(g2260B),.A2(I5297B),.A1(I5296B));
NAND4_X1 U_g7986B (.ZN(g7986B),.A4(g7550B),.A3(g2172B),.A2(FE_OFN80_g2175B),.A1(FE_OFN88_g2178B));
NAND2_X1 U_g5226B (.ZN(g5226B),.A2(I8671B),.A1(I8670B));
NAND2_X1 U_g8512B (.ZN(g8512B),.A2(g8366B),.A1(g3723B));
NAND2_X1 U_I16046B (.ZN(I16046B),.A2(I16044B),.A1(g10432B));
NAND2_X1 U_I13504B (.ZN(I13504B),.A2(g8247B),.A1(g677B));
NAND2_X1 U_g10447B (.ZN(g10447B),.A2(g5360B),.A1(g10363B));
NAND2_X1 U_g2167B (.ZN(g2167B),.A2(I5106B),.A1(I5105B));
NAND2_X1 U_I8804B (.ZN(I8804B),.A2(I8803B),.A1(g4677B));
NAND2_X1 U_g10472B (.ZN(g10472B),.A2(I16017B),.A1(I16016B));
NAND2_X1 U_I17487B (.ZN(I17487B),.A2(I17485B),.A1(g11474B));
NAND2_X1 U_I4995B (.ZN(I4995B),.A2(g309B),.A1(g416B));
NAND2_X1 U_I12093B (.ZN(I12093B),.A2(I12092B),.A1(g5810B));
NAND4_X1 U_g7987B (.ZN(g7987B),.A4(FE_OFN96_g2169B),.A3(g7562B),.A2(FE_OFN80_g2175B),.A1(FE_OFN88_g2178B));
NAND2_X1 U_g5227B (.ZN(g5227B),.A2(I8678B),.A1(I8677B));
NAND2_X1 U_I5126B (.ZN(I5126B),.A2(g1389B),.A1(g1386B));
NAND2_X1 U_g2321B (.ZN(g2321B),.A2(I5373B),.A1(I5372B));
NAND2_X1 U_g7547B (.ZN(g7547B),.A2(I11975B),.A1(I11974B));
NAND2_X1 U_I17306B (.ZN(I17306B),.A2(I17305B),.A1(g11232B));
NAND3_X1 U_g6548B (.ZN(g6548B),.A3(g6122B),.A2(g6124B),.A1(g826B));
NAND2_X1 U_I11995B (.ZN(I11995B),.A2(g127B),.A1(g6035B));
NAND2_X1 U_I7225B (.ZN(I7225B),.A2(I7223B),.A1(g1781B));
NAND2_X1 U_I11261B (.ZN(I11261B),.A2(g826B),.A1(g6775B));
NAND3_X1 U_g8843B (.ZN(g8843B),.A3(g8545B),.A2(g8757B),.A1(g8542B));
NAND2_X1 U_g2938B (.ZN(g2938B),.A2(I6111B),.A1(I6110B));
NAND2_X1 U_I4942B (.ZN(I4942B),.A2(I4941B),.A1(g396B));
NAND2_X1 U_g10394B (.ZN(g10394B),.A2(I15900B),.A1(I15899B));
NAND2_X1 U_g8549B (.ZN(g8549B),.A2(g8390B),.A1(g5527B));
NAND2_X1 U_g3070B (.ZN(g3070B),.A2(g1206B),.A1(g2016B));
NAND2_X1 U_I4954B (.ZN(I4954B),.A2(g327B),.A1(g401B));
NAND2_X1 U_I5023B (.ZN(I5023B),.A2(g1275B),.A1(g995B));
NAND2_X1 U_g10446B (.ZN(g10446B),.A2(g5350B),.A1(g10438B));
NAND2_X1 U_I16081B (.ZN(I16081B),.A2(I16079B),.A1(g10363B));
NAND2_X1 U_I8641B (.ZN(I8641B),.A2(I8640B),.A1(g4278B));
NAND2_X1 U_I6178B (.ZN(I6178B),.A2(I6176B),.A1(g197B));
NAND2_X1 U_I12075B (.ZN(I12075B),.A2(I12074B),.A1(g6015B));
NAND2_X1 U_I5127B (.ZN(I5127B),.A2(I5126B),.A1(g1386B));
NAND2_X1 U_I5451B (.ZN(I5451B),.A2(I5449B),.A1(g991B));
NAND2_X1 U_g4168B (.ZN(g4168B),.A2(I7323B),.A1(I7322B));
NAND2_X1 U_I6288B (.ZN(I6288B),.A2(I6287B),.A1(g2091B));
NAND2_X1 U_I8179B (.ZN(I8179B),.A2(I8178B),.A1(g3685B));
NAND2_X1 U_I4912B (.ZN(I4912B),.A2(I4910B),.A1(g318B));
NAND2_X1 U_I6805B (.ZN(I6805B),.A2(g471B),.A1(g3268B));
NAND3_X1 U_g3766B (.ZN(g3766B),.A3(g2493B),.A2(g3222B),.A1(g2439B));
NAND2_X1 U_g3087B (.ZN(g3087B),.A2(I6289B),.A1(I6288B));
NAND2_X1 U_I17486B (.ZN(I17486B),.A2(I17485B),.A1(g11233B));
NAND2_X1 U_I4929B (.ZN(I4929B),.A2(I4928B),.A1(g391B));
NAND2_X1 U_I15890B (.ZN(I15890B),.A2(g10285B),.A1(g853B));
NAND2_X1 U_I16331B (.ZN(I16331B),.A2(I16330B),.A1(g10387B));
NAND2_X1 U_I9575B (.ZN(I9575B),.A2(I9574B),.A1(g5608B));
NAND2_X1 U_I13887B (.ZN(I13887B),.A2(I13886B),.A1(g8267B));
NAND2_X1 U_g5308B (.ZN(g5308B),.A2(I8788B),.A1(I8787B));
NAND2_X1 U_I13529B (.ZN(I13529B),.A2(g8253B),.A1(g704B));
NAND2_X1 U_I6208B (.ZN(I6208B),.A2(I6207B),.A1(g5188B));
NAND2_X1 U_g5217B (.ZN(g5217B),.A2(I8642B),.A1(I8641B));
NAND2_X1 U_I5316B (.ZN(I5316B),.A2(I5315B),.A1(g1032B));
NAND2_X1 U_g2111B (.ZN(g2111B),.A2(I5007B),.A1(I5006B));
NAND2_X1 U_g10366B (.ZN(g10366B),.A2(g5392B),.A1(g10285B));
NAND2_X1 U_I5034B (.ZN(I5034B),.A2(g1019B),.A1(g1015B));
NAND2_X1 U_I13869B (.ZN(I13869B),.A2(I13867B),.A1(g1403B));
NAND2_X1 U_I13868B (.ZN(I13868B),.A2(I13867B),.A1(g8264B));
NAND2_X1 U_I15999B (.ZN(I15999B),.A2(FE_OFN247_g1771B),.A1(g10432B));
NAND2_X1 U_I13259B (.ZN(I13259B),.A2(I13258B),.A1(g1900B));
NAND4_X1 U_g3261B (.ZN(g3261B),.A4(g2202B),.A3(g2211B),.A2(g2222B),.A1(g2229B));
NAND2_X1 U_g10481B (.ZN(g10481B),.A2(I16074B),.A1(I16073B));
NAND2_X1 U_g2180B (.ZN(g2180B),.A2(I5137B),.A1(I5136B));
NAND3_X1 U_g4976B (.ZN(g4976B),.A3(g3807B),.A2(g4604B),.A1(g2310B));
NAND2_X1 U_g8506B (.ZN(g8506B),.A2(g8366B),.A1(g3475B));
NAND2_X1 U_g2380B (.ZN(g2380B),.A2(I5461B),.A1(I5460B));
NAND2_X1 U_I13258B (.ZN(I13258B),.A2(g8153B),.A1(g1900B));
NAND2_X1 U_I5013B (.ZN(I5013B),.A2(g1011B),.A1(g1007B));
NAND2_X1 U_g5196B (.ZN(g5196B),.A2(I8606B),.A1(I8605B));
NAND2_X1 U_I10930B (.ZN(I10930B),.A2(g5555B),.A1(g5863B));
NAND2_X1 U_I6770B (.ZN(I6770B),.A2(g382B),.A1(g3257B));
NAND2_X1 U_g11449B (.ZN(g11449B),.A2(I17402B),.A1(I17401B));
NAND2_X1 U_g11448B (.ZN(g11448B),.A2(I17395B),.A1(I17394B));
NAND2_X1 U_I15717B (.ZN(I15717B),.A2(I15716B),.A1(g10231B));
NAND2_X1 U_I5317B (.ZN(I5317B),.A2(I5315B),.A1(g1027B));
NAND2_X1 U_I14210B (.ZN(I14210B),.A2(I14209B),.A1(g8824B));
NAND2_X1 U_I17569B (.ZN(I17569B),.A2(I17567B),.A1(g1610B));
NAND2_X1 U_I13878B (.ZN(I13878B),.A2(I13876B),.A1(g1444B));
NAND2_X1 U_g8545B (.ZN(g8545B),.A2(g8390B),.A1(g3710B));
NAND2_X1 U_g2515B (.ZN(g2515B),.A2(I5606B),.A1(I5605B));
NAND2_X1 U_I14443B (.ZN(I14443B),.A2(I14442B),.A1(g8970B));
NAND2_X1 U_g7557B (.ZN(g7557B),.A2(I11997B),.A1(I11996B));
NAND2_X1 U_g8180B (.ZN(g8180B),.A2(I13091B),.A1(I13090B));
NAND2_X1 U_I14279B (.ZN(I14279B),.A2(I14277B),.A1(g1828B));
NAND2_X1 U_I17568B (.ZN(I17568B),.A2(I17567B),.A1(g11496B));
NAND2_X1 U_I13886B (.ZN(I13886B),.A2(g1440B),.A1(g8267B));
NAND2_X1 U_I7322B (.ZN(I7322B),.A2(I7321B),.A1(g3047B));
NAND2_X1 U_I6990B (.ZN(I6990B),.A2(I6988B),.A1(g986B));
NAND2_X1 U_I14278B (.ZN(I14278B),.A2(I14277B),.A1(g8847B));
NAND2_X1 U_I7033B (.ZN(I7033B),.A2(g1868B),.A1(g3089B));
NAND2_X1 U_I9006B (.ZN(I9006B),.A2(FE_OFN252_g1791B),.A1(g4492B));
NAND2_X1 U_g8507B (.ZN(g8507B),.A2(g8366B),.A1(g3738B));
NAND2_X1 U_I5460B (.ZN(I5460B),.A2(I5459B),.A1(g1240B));
NAND2_X1 U_g4588B (.ZN(g4588B),.A2(FE_OFN325_g18B),.A1(g3440B));
NAND2_X1 U_I4986B (.ZN(I4986B),.A2(I4985B),.A1(g999B));
NAND3_X1 U_g3247B (.ZN(g3247B),.A3(g2571B),.A2(g2564B),.A1(g1828B));
NAND2_X1 U_I8651B (.ZN(I8651B),.A2(I8650B),.A1(g4824B));
NAND2_X1 U_I13545B (.ZN(I13545B),.A2(I13544B),.A1(g713B));
NAND2_X1 U_g8628B (.ZN(g8628B),.A2(I13895B),.A1(I13894B));
NAND2_X1 U_I6138B (.ZN(I6138B),.A2(I6136B),.A1(g378B));
NAND2_X1 U_I12074B (.ZN(I12074B),.A2(g174B),.A1(g6015B));
NAND2_X1 U_g8630B (.ZN(g8630B),.A2(I13909B),.A1(I13908B));
NAND2_X1 U_I13078B (.ZN(I13078B),.A2(I13076B),.A1(g7963B));
NAND2_X1 U_I6109B (.ZN(I6109B),.A2(g1494B),.A1(g2205B));
NAND2_X1 U_g8300B (.ZN(g8300B),.A2(I13260B),.A1(I13259B));
NAND2_X1 U_I5501B (.ZN(I5501B),.A2(I5500B),.A1(g1255B));
NAND2_X1 U_I17586B (.ZN(I17586B),.A2(I17584B),.A1(g11515B));
NAND2_X1 U_I12092B (.ZN(I12092B),.A2(g1490B),.A1(g5810B));
NAND2_X1 U_I13901B (.ZN(I13901B),.A2(I13900B),.A1(g8261B));
NAND2_X1 U_I8795B (.ZN(I8795B),.A2(g1145B),.A1(g4672B));
NAND2_X1 U_I6201B (.ZN(I6201B),.A2(I6199B),.A1(g766B));
NAND2_X1 U_I14217B (.ZN(I14217B),.A2(I14216B),.A1(g8826B));
NAND2_X1 U_I9007B (.ZN(I9007B),.A2(I9006B),.A1(g4492B));
NAND2_X1 U_I13561B (.ZN(I13561B),.A2(I13559B),.A1(g8263B));
NAND2_X1 U_I15716B (.ZN(I15716B),.A2(g10229B),.A1(g10231B));
NAND2_X1 U_I6449B (.ZN(I6449B),.A2(I6447B),.A1(FE_OFN236_g1776B));
NAND2_X1 U_I13295B (.ZN(I13295B),.A2(I13293B),.A1(g8161B));
NAND2_X1 U_I4987B (.ZN(I4987B),.A2(I4985B),.A1(g1003B));
NAND2_X1 U_I6715B (.ZN(I6715B),.A2(I6714B),.A1(g2961B));
NAND2_X1 U_I17493B (.ZN(I17493B),.A2(I17492B),.A1(g11430B));
NAND2_X1 U_I12215B (.ZN(I12215B),.A2(I12214B),.A1(g7061B));
NAND2_X1 U_g2372B (.ZN(g2372B),.A2(I5451B),.A1(I5450B));
NAND2_X1 U_g7062B (.ZN(g7062B),.A2(I11263B),.A1(I11262B));
NAND2_X1 U_g2988B (.ZN(g2988B),.A2(I6226B),.A1(I6225B));
NAND2_X1 U_I13309B (.ZN(I13309B),.A2(I13307B),.A1(g617B));
NAND2_X1 U_g8839B (.ZN(g8839B),.A2(FE_OFN223_g4401B),.A1(g8603B));
NAND2_X1 U_g2555B (.ZN(g2555B),.A2(I5677B),.A1(I5676B));
NAND2_X1 U_g3662B (.ZN(g3662B),.A2(I6827B),.A1(I6826B));
NAND2_X1 U_I13308B (.ZN(I13308B),.A2(I13307B),.A1(g8190B));
NAND2_X1 U_g2792B (.ZN(g2792B),.A2(I5880B),.A1(I5879B));
NAND2_X1 U_g4117B (.ZN(g4117B),.A2(g3061B),.A1(g3041B));
NAND2_X1 U_I8543B (.ZN(I8543B),.A2(g486B),.A1(g4218B));
NAND2_X1 U_g11549B (.ZN(g11549B),.A2(I17586B),.A1(I17585B));
NAND2_X1 U_I6881B (.ZN(I6881B),.A2(I6879B),.A1(g1351B));
NAND2_X1 U_I12138B (.ZN(I12138B),.A2(I12136B),.A1(g131B));
NAND2_X1 U_I8729B (.ZN(I8729B),.A2(I8728B),.A1(g4605B));
NAND2_X1 U_I14216B (.ZN(I14216B),.A2(g605B),.A1(g8826B));
NAND2_X1 U_g10384B (.ZN(g10384B),.A2(I15872B),.A1(I15871B));
NAND2_X1 U_I13260B (.ZN(I13260B),.A2(I13258B),.A1(g8153B));
NAND2_X1 U_g2776B (.ZN(g2776B),.A2(I5867B),.A1(I5866B));
NAND2_X1 U_I8513B (.ZN(I8513B),.A2(g3513B),.A1(g4873B));
NAND2_X1 U_I13559B (.ZN(I13559B),.A2(g8263B),.A1(g722B));
NAND2_X1 U_I8178B (.ZN(I8178B),.A2(FE_OFN253_g1786B),.A1(g3685B));
NAND2_X1 U_g3631B (.ZN(g3631B),.A2(I6794B),.A1(I6793B));
NAND2_X1 U_I6487B (.ZN(I6487B),.A2(g1227B),.A1(g2306B));
NAND2_X1 U_I16080B (.ZN(I16080B),.A2(I16079B),.A1(g849B));
NAND2_X1 U_I13893B (.ZN(I13893B),.A2(g1436B),.A1(g8266B));
NAND2_X1 U_I12115B (.ZN(I12115B),.A2(I12113B),.A1(g162B));
NAND2_X1 U_I6748B (.ZN(I6748B),.A2(I6746B),.A1(g1453B));
NAND2_X1 U_I13544B (.ZN(I13544B),.A2(g8259B),.A1(g713B));
NAND2_X1 U_I5484B (.ZN(I5484B),.A2(g1011B),.A1(g1250B));
NAND2_X1 U_I4928B (.ZN(I4928B),.A2(g321B),.A1(g391B));
NAND2_X1 U_I6226B (.ZN(I6226B),.A2(I6224B),.A1(g1346B));
NAND2_X1 U_I8805B (.ZN(I8805B),.A2(I8803B),.A1(g1113B));
NAND2_X1 U_I4930B (.ZN(I4930B),.A2(I4928B),.A1(g321B));
NAND2_X1 U_I15880B (.ZN(I15880B),.A2(I15878B),.A1(FE_OFN251_g1801B));
NAND2_X1 U_I14265B (.ZN(I14265B),.A2(I14263B),.A1(g1814B));
NAND2_X1 U_I16031B (.ZN(I16031B),.A2(I16030B),.A1(g829B));
NAND2_X1 U_g3585B (.ZN(g3585B),.A2(I6748B),.A1(I6747B));
NAND4_X1 U_g3041B (.ZN(g3041B),.A4(g2382B),.A3(g2374B),.A2(g2399B),.A1(g2364B));
NAND2_X1 U_g8933B (.ZN(g8933B),.A2(I14272B),.A1(I14271B));
NAND2_X1 U_I16330B (.ZN(I16330B),.A2(g4997B),.A1(g10387B));
NAND2_X1 U_I13267B (.ZN(I13267B),.A2(I13265B),.A1(g8154B));
NAND2_X1 U_I13294B (.ZN(I13294B),.A2(I13293B),.A1(g1882B));
NAND2_X1 U_g10231B (.ZN(g10231B),.A2(I15617B),.A1(I15616B));
NAND2_X1 U_I14442B (.ZN(I14442B),.A2(g1834B),.A1(g8970B));
NAND2_X1 U_I6793B (.ZN(I6793B),.A2(I6792B),.A1(g2959B));
NAND2_X1 U_I4966B (.ZN(I4966B),.A2(I4964B),.A1(g330B));
NAND2_X1 U_I8752B (.ZN(I8752B),.A2(I8750B),.A1(g1125B));
NAND2_X1 U_I15432B (.ZN(I15432B),.A2(I15430B),.A1(g9995B));
NAND2_X1 U_I12214B (.ZN(I12214B),.A2(g2518B),.A1(g7061B));
NAND2_X1 U_g10511B (.ZN(g10511B),.A2(g6032B),.A1(g10438B));
NAND2_X1 U_g3011B (.ZN(g3011B),.A2(g2382B),.A1(g591B));
NAND2_X1 U_g5103B (.ZN(g5103B),.A2(I8481B),.A1(I8480B));
NAND2_X1 U_I16087B (.ZN(I16087B),.A2(I16086B),.A1(g861B));
NAND2_X1 U_g3734B (.ZN(g3734B),.A2(g599B),.A1(g3039B));
NAND2_X1 U_I6664B (.ZN(I6664B),.A2(g2776B),.A1(g2792B));
NAND2_X1 U_g8882B (.ZN(g8882B),.A2(I14218B),.A1(I14217B));
NAND2_X1 U_I4955B (.ZN(I4955B),.A2(I4954B),.A1(g401B));
NAND2_X1 U_I8786B (.ZN(I8786B),.A2(g1141B),.A1(g4639B));
NAND3_X1 U_g3992B (.ZN(g3992B),.A3(g2990B),.A2(g2550B),.A1(g2571B));
NAND2_X1 U_g10480B (.ZN(g10480B),.A2(I16067B),.A1(I16066B));
NAND2_X1 U_I11915B (.ZN(I11915B),.A2(I11914B),.A1(g5803B));
NAND2_X1 U_I8770B (.ZN(I8770B),.A2(g1133B),.A1(g4619B));
NAND2_X1 U_I5516B (.ZN(I5516B),.A2(g1019B),.A1(g1260B));
NAND2_X1 U_g8541B (.ZN(g8541B),.A2(g8390B),.A1(g4001B));
NAND2_X1 U_I6188B (.ZN(I6188B),.A2(I6186B),.A1(g466B));
NAND2_X1 U_g5147B (.ZN(g5147B),.A2(I8545B),.A1(I8544B));
NAND3_X1 U_g8744B (.ZN(g8744B),.A3(I9273B),.A2(g46B),.A1(g8617B));
NAND2_X1 U_I5892B (.ZN(I5892B),.A2(I5891B),.A1(g750B));
NAND2_X1 U_g8558B (.ZN(g8558B),.A2(I13767B),.A1(I13766B));
NAND2_X1 U_I15258B (.ZN(I15258B),.A2(I15256B),.A1(g9968B));
NAND2_X1 U_I13266B (.ZN(I13266B),.A2(I13265B),.A1(g1909B));
NAND2_X1 U_I8787B (.ZN(I8787B),.A2(I8786B),.A1(g4639B));
NAND2_X1 U_I6826B (.ZN(I6826B),.A2(I6825B),.A1(g3281B));
NAND2_X1 U_I17283B (.ZN(I17283B),.A2(I17281B),.A1(g11219B));
NAND3_X1 U_g5013B (.ZN(g5013B),.A3(g3205B),.A2(g3247B),.A1(g4749B));
NAND2_X1 U_I17492B (.ZN(I17492B),.A2(g3623B),.A1(g11430B));
NAND2_X1 U_g8511B (.ZN(g8511B),.A2(g8366B),.A1(g5277B));
NAND2_X1 U_I16079B (.ZN(I16079B),.A2(g10363B),.A1(g849B));
NAND2_X1 U_I5035B (.ZN(I5035B),.A2(I5034B),.A1(g1015B));
NAND2_X1 U_I5517B (.ZN(I5517B),.A2(I5516B),.A1(g1260B));
NAND2_X1 U_I7223B (.ZN(I7223B),.A2(g1781B),.A1(g2981B));
NAND2_X1 U_I16086B (.ZN(I16086B),.A2(g10430B),.A1(g861B));
NAND2_X1 U_g5317B (.ZN(g5317B),.A2(I8797B),.A1(I8796B));
NAND2_X1 U_I15879B (.ZN(I15879B),.A2(I15878B),.A1(g10359B));
NAND2_X1 U_I15878B (.ZN(I15878B),.A2(FE_OFN251_g1801B),.A1(g10359B));
NAND2_X1 U_I12114B (.ZN(I12114B),.A2(I12113B),.A1(g6002B));
NAND2_X1 U_I12107B (.ZN(I12107B),.A2(I12106B),.A1(g6042B));
NAND2_X1 U_g2500B (.ZN(g2500B),.A2(g182B),.A1(g178B));
NAND2_X1 U_I15994B (.ZN(I15994B),.A2(I15992B),.A1(g2677B));
NAND4_X1 U_g7934B (.ZN(g7934B),.A4(g7550B),.A3(FE_OFN91_g2172B),.A2(FE_OFN80_g2175B),.A1(g6941B));
NAND2_X1 U_g10469B (.ZN(g10469B),.A2(g5999B),.A1(g10430B));
NAND2_X1 U_I14264B (.ZN(I14264B),.A2(I14263B),.A1(g8843B));
NAND2_X1 U_I6448B (.ZN(I6448B),.A2(I6447B),.A1(g2264B));
NAND2_X1 U_I13285B (.ZN(I13285B),.A2(I13283B),.A1(g8159B));
NAND2_X1 U_g10468B (.ZN(g10468B),.A2(I16001B),.A1(I16000B));
NAND2_X1 U_I6827B (.ZN(I6827B),.A2(I6825B),.A1(g770B));
NAND2_X1 U_g8623B (.ZN(g8623B),.A2(I13878B),.A1(I13877B));
NAND2_X1 U_I13900B (.ZN(I13900B),.A2(g1428B),.A1(g8261B));
NAND2_X1 U_g2795B (.ZN(g2795B),.A2(I5893B),.A1(I5892B));
NAND2_X1 U_I8575B (.ZN(I8575B),.A2(g496B),.A1(g4234B));
NAND2_X1 U_I14209B (.ZN(I14209B),.A2(g599B),.A1(g8824B));
NAND2_X1 U_I13560B (.ZN(I13560B),.A2(I13559B),.A1(g722B));
NAND2_X1 U_I8715B (.ZN(I8715B),.A2(g4052B),.A1(g4601B));
NAND2_X1 U_I8604B (.ZN(I8604B),.A2(g506B),.A1(g4259B));
NAND2_X1 U_I16017B (.ZN(I16017B),.A2(I16015B),.A1(g1781B));
NAND2_X1 U_I4941B (.ZN(I4941B),.A2(g324B),.A1(g396B));
NAND2_X1 U_g2205B (.ZN(g2205B),.A2(I5166B),.A1(I5165B));
NAND3_X1 U_g3753B (.ZN(g3753B),.A3(g2800B),.A2(g2364B),.A1(g2382B));
NAND2_X1 U_I6467B (.ZN(I6467B),.A2(g2479B),.A1(g23B));
NAND2_X1 U_I14614B (.ZN(I14614B),.A2(I14612B),.A1(g611B));
NAND2_X1 U_g2104B (.ZN(g2104B),.A2(I4966B),.A1(I4965B));
NAND2_X1 U_g2099B (.ZN(g2099B),.A2(I4943B),.A1(I4942B));
NAND2_X1 U_I16023B (.ZN(I16023B),.A2(FE_OFN253_g1786B),.A1(g10438B));
NAND2_X1 U_g10479B (.ZN(g10479B),.A2(I16060B),.A1(I16059B));
NAND3_X1 U_g8737B (.ZN(g8737B),.A3(g8688B),.A2(FE_OFN200_g4921B),.A1(g1975B));
NAND2_X1 U_g5942B (.ZN(g5942B),.A2(I9576B),.A1(I9575B));
NAND2_X1 U_g10478B (.ZN(g10478B),.A2(I16053B),.A1(I16052B));
NAND2_X1 U_I12004B (.ZN(I12004B),.A2(I12002B),.A1(g153B));
NAND2_X1 U_I4911B (.ZN(I4911B),.A2(I4910B),.A1(g386B));
NAND2_X1 U_I11914B (.ZN(I11914B),.A2(g1494B),.A1(g5803B));
NAND2_X1 U_g7960B (.ZN(g7960B),.A2(g5573B),.A1(g7409B));
NAND2_X1 U_I5295B (.ZN(I5295B),.A2(g798B),.A1(g794B));
NAND2_X1 U_I12106B (.ZN(I12106B),.A2(g135B),.A1(g6042B));
NAND2_X1 U_I8728B (.ZN(I8728B),.A2(g1117B),.A1(g4605B));
NAND2_X1 U_g3681B (.ZN(g3681B),.A2(I6838B),.A1(I6837B));
NAND2_X1 U_I11907B (.ZN(I11907B),.A2(g1474B),.A1(g5838B));
NAND2_X1 U_I13907B (.ZN(I13907B),.A2(g1432B),.A1(g8265B));
NAND2_X1 U_I8730B (.ZN(I8730B),.A2(I8728B),.A1(g1117B));
NAND2_X1 U_g8551B (.ZN(g8551B),.A2(g8390B),.A1(g3967B));
NAND2_X1 U_I4980B (.ZN(I4980B),.A2(I4978B),.A1(g333B));
NAND2_X1 U_g2961B (.ZN(g2961B),.A2(I6178B),.A1(I6177B));
NAND2_X1 U_g6019B (.ZN(g6019B),.A2(FE_OFN200_g4921B),.A1(g617B));
NAND2_X1 U_I16016B (.ZN(I16016B),.A2(I16015B),.A1(g10441B));
NAND2_X1 U_I11935B (.ZN(I11935B),.A2(g1458B),.A1(g5857B));
NAND2_X1 U_I8678B (.ZN(I8678B),.A2(I8676B),.A1(g1027B));
NAND2_X1 U_I17051B (.ZN(I17051B),.A2(g11249B),.A1(g10923B));
NAND2_X1 U_g4482B (.ZN(g4482B),.A2(I7865B),.A1(I7864B));
NAND2_X1 U_g7592B (.ZN(g7592B),.A2(I12108B),.A1(I12107B));
NAND2_X1 U_g3460B (.ZN(g3460B),.A2(I6666B),.A1(I6665B));
NAND4_X1 U_g7932B (.ZN(g7932B),.A4(FE_OFN96_g2169B),.A3(FE_OFN91_g2172B),.A2(FE_OFN80_g2175B),.A1(g6941B));
NAND2_X1 U_g7624B (.ZN(g7624B),.A2(I12216B),.A1(I12215B));
NAND4_X1 U_g7953B (.ZN(g7953B),.A4(g7550B),.A3(g7562B),.A2(g7574B),.A1(g6941B));
NAND2_X1 U_g8414B (.ZN(g8414B),.A2(I13554B),.A1(I13553B));
NAND2_X1 U_I6168B (.ZN(I6168B),.A2(I6166B),.A1(g153B));
NAND2_X1 U_I5229B (.ZN(I5229B),.A2(g148B),.A1(g182B));
NAND2_X1 U_I6772B (.ZN(I6772B),.A2(I6770B),.A1(g382B));
NAND2_X1 U_I16030B (.ZN(I16030B),.A2(g10430B),.A1(g829B));
NAND2_X1 U_I13284B (.ZN(I13284B),.A2(I13283B),.A1(g1927B));
NAND2_X1 U_I16065B (.ZN(I16065B),.A2(FE_OFN237_g1806B),.A1(g10428B));
NAND2_X1 U_g2947B (.ZN(g2947B),.A2(I6138B),.A1(I6137B));
NAND2_X1 U_I7321B (.ZN(I7321B),.A2(g1231B),.A1(g3047B));
NAND2_X1 U_g2437B (.ZN(g2437B),.A2(I5530B),.A1(I5529B));
NAND2_X1 U_g2102B (.ZN(g2102B),.A2(I4956B),.A1(I4955B));
NAND2_X1 U_I17282B (.ZN(I17282B),.A2(I17281B),.A1(g11221B));
NAND2_X1 U_I5620B (.ZN(I5620B),.A2(I5618B),.A1(FE_OFN247_g1771B));
NAND2_X1 U_I8664B (.ZN(I8664B),.A2(I8662B),.A1(g476B));
NAND2_X1 U_g7524B (.ZN(g7524B),.A2(I11916B),.A1(I11915B));
NAND2_X1 U_g7717B (.ZN(g7717B),.A2(g1950B),.A1(g6863B));
NAND2_X1 U_I16467B (.ZN(I16467B),.A2(g10518B),.A1(g10716B));
NAND2_X1 U_I4972B (.ZN(I4972B),.A2(I4971B),.A1(g991B));
NAND2_X1 U_I13554B (.ZN(I13554B),.A2(I13552B),.A1(g8262B));
NAND2_X1 U_I16037B (.ZN(I16037B),.A2(FE_OFN252_g1791B),.A1(g10363B));
NAND2_X1 U_g8302B (.ZN(g8302B),.A2(I13274B),.A1(I13273B));
NAND2_X1 U_I4943B (.ZN(I4943B),.A2(I4941B),.A1(g324B));
NAND2_X1 U_I5485B (.ZN(I5485B),.A2(I5484B),.A1(g1250B));
NAND2_X1 U_g5527B (.ZN(g5527B),.A2(g4749B),.A1(g3978B));
NAND2_X1 U_I10509B (.ZN(I10509B),.A2(I10507B),.A1(g786B));
NAND2_X1 U_g7599B (.ZN(g7599B),.A2(I12145B),.A1(I12144B));
NAND2_X1 U_I10508B (.ZN(I10508B),.A2(I10507B),.A1(g6221B));
NAND2_X1 U_I6126B (.ZN(I6126B),.A2(I6124B),.A1(g1419B));
NAND2_X1 U_I8671B (.ZN(I8671B),.A2(I8669B),.A1(g814B));
NAND2_X1 U_I6760B (.ZN(I6760B),.A2(g1448B),.A1(g2943B));
NAND2_X1 U_g3626B (.ZN(g3626B),.A2(I6779B),.A1(I6778B));
NAND2_X1 U_I11973B (.ZN(I11973B),.A2(g1462B),.A1(g5852B));
NAND2_X1 U_g2389B (.ZN(g2389B),.A2(I5470B),.A1(I5469B));
NAND2_X1 U_I15617B (.ZN(I15617B),.A2(I15615B),.A1(g10153B));
NAND2_X1 U_g5277B (.ZN(g5277B),.A2(g4538B),.A1(g3734B));
NAND2_X1 U_I5005B (.ZN(I5005B),.A2(g312B),.A1(g421B));
NAND2_X1 U_I6779B (.ZN(I6779B),.A2(I6777B),.A1(g650B));
NAND2_X1 U_I6665B (.ZN(I6665B),.A2(I6664B),.A1(g2792B));
NAND2_X1 U_I8589B (.ZN(I8589B),.A2(g501B),.A1(g4251B));
NAND2_X1 U_g8412B (.ZN(g8412B),.A2(I13546B),.A1(I13545B));
NAND2_X1 U_g2963B (.ZN(g2963B),.A2(I6188B),.A1(I6187B));
NAND2_X1 U_I12045B (.ZN(I12045B),.A2(g1486B),.A1(g5814B));
NAND2_X1 U_I16053B (.ZN(I16053B),.A2(I16051B),.A1(g10434B));
NAND2_X1 U_g2109B (.ZN(g2109B),.A2(I4997B),.A1(I4996B));
NAND2_X1 U_g11418B (.ZN(g11418B),.A2(I17307B),.A1(I17306B));
NAND2_X1 U_I13539B (.ZN(I13539B),.A2(I13537B),.A1(g8157B));
NAND2_X1 U_g10475B (.ZN(g10475B),.A2(I16032B),.A1(I16031B));
NAND2_X1 U_I5324B (.ZN(I5324B),.A2(I5323B),.A1(g1336B));
NAND2_X1 U_I13538B (.ZN(I13538B),.A2(I13537B),.A1(g658B));
NAND2_X1 U_I5469B (.ZN(I5469B),.A2(I5468B),.A1(g1245B));
NAND2_X1 U_I5540B (.ZN(I5540B),.A2(I5538B),.A1(g1023B));
NAND2_X1 U_I17505B (.ZN(I17505B),.A2(I17503B),.A1(g5269B));
NAND2_X1 U_I11241B (.ZN(I11241B),.A2(g790B),.A1(g6760B));
NAND2_X1 U_I8803B (.ZN(I8803B),.A2(g1113B),.A1(g4677B));
NAND2_X1 U_I12061B (.ZN(I12061B),.A2(I12060B),.A1(g5824B));
NAND2_X1 U_I8780B (.ZN(I8780B),.A2(I8778B),.A1(g1137B));
NAND3_X1 U_g8745B (.ZN(g8745B),.A3(I9265B),.A2(g47B),.A1(g8617B));
NAND2_X1 U_I4979B (.ZN(I4979B),.A2(I4978B),.A1(g411B));
NAND2_X1 U_g8109B (.ZN(g8109B),.A2(I11360B),.A1(g48B));
NAND2_X1 U_g8309B (.ZN(g8309B),.A2(I13309B),.A1(I13308B));
NAND2_X1 U_g6758B (.ZN(g6758B),.A2(I10771B),.A1(I10770B));
NAND2_X1 U_I16009B (.ZN(I16009B),.A2(I16007B),.A1(FE_OFN236_g1776B));
NAND2_X1 U_I15616B (.ZN(I15616B),.A2(I15615B),.A1(g10043B));
NAND2_X1 U_I8662B (.ZN(I8662B),.A2(g476B),.A1(g4286B));
NAND2_X1 U_I16008B (.ZN(I16008B),.A2(I16007B),.A1(g10434B));
NAND2_X1 U_I13515B (.ZN(I13515B),.A2(I13513B),.A1(g8248B));
NAND2_X1 U_I13991B (.ZN(I13991B),.A2(I13990B),.A1(g622B));
NAND2_X1 U_g11276B (.ZN(g11276B),.A2(I17053B),.A1(I17052B));
NAND2_X1 U_I15900B (.ZN(I15900B),.A2(I15898B),.A1(g10359B));
NAND2_X1 U_g2419B (.ZN(g2419B),.A2(I5502B),.A1(I5501B));
NAND2_X1 U_I16074B (.ZN(I16074B),.A2(I16072B),.A1(g10438B));
NAND2_X1 U_I10769B (.ZN(I10769B),.A2(FE_OFN251_g1801B),.A1(g5944B));
NAND2_X1 U_I7323B (.ZN(I7323B),.A2(I7321B),.A1(g1231B));
NAND2_X1 U_g7978B (.ZN(g7978B),.A2(g736B),.A1(g7697B));
NAND2_X1 U_I7875B (.ZN(I7875B),.A2(g810B),.A1(g4109B));
NAND2_X1 U_I8562B (.ZN(I8562B),.A2(I8561B),.A1(g4227B));
NAND2_X1 U_I15892B (.ZN(I15892B),.A2(I15890B),.A1(g10285B));
NAND2_X1 U_g3771B (.ZN(g3771B),.A2(I6990B),.A1(I6989B));
NAND2_X1 U_I8605B (.ZN(I8605B),.A2(I8604B),.A1(g4259B));
NAND2_X1 U_g10153B (.ZN(g10153B),.A2(I15453B),.A1(I15452B));
NAND2_X1 U_g5295B (.ZN(g5295B),.A2(I8763B),.A1(I8762B));
NAND2_X1 U_I8751B (.ZN(I8751B),.A2(I8750B),.A1(g4613B));
NAND2_X1 U_I15907B (.ZN(I15907B),.A2(I15906B),.A1(g6899B));
NAND2_X1 U_I5136B (.ZN(I5136B),.A2(I5135B),.A1(g521B));
NAND2_X1 U_I11263B (.ZN(I11263B),.A2(I11261B),.A1(g826B));
NAND2_X1 U_I14204B (.ZN(I14204B),.A2(I14202B),.A1(g591B));
NAND2_X1 U_g8881B (.ZN(g8881B),.A2(I14211B),.A1(I14210B));
NAND2_X1 U_g2105B (.ZN(g2105B),.A2(I4973B),.A1(I4972B));
NAND3_X1 U_g5557B (.ZN(g5557B),.A3(g3011B),.A2(g3071B),.A1(g4538B));
NAND2_X1 U_I5230B (.ZN(I5230B),.A2(I5229B),.A1(g182B));
NAND2_X1 U_I8669B (.ZN(I8669B),.A2(g814B),.A1(g4831B));
NAND2_X1 U_g10474B (.ZN(g10474B),.A2(I16025B),.A1(I16024B));
NAND2_X1 U_I8772B (.ZN(I8772B),.A2(I8770B),.A1(g1133B));
NAND2_X1 U_g2445B (.ZN(g2445B),.A2(I5540B),.A1(I5539B));
NAND2_X1 U_g8006B (.ZN(g8006B),.A2(g7717B),.A1(g5552B));
NAND2_X1 U_I10932B (.ZN(I10932B),.A2(I10930B),.A1(g5555B));
NAND2_X1 U_I17504B (.ZN(I17504B),.A2(I17503B),.A1(g11430B));
NAND2_X1 U_I5137B (.ZN(I5137B),.A2(I5135B),.A1(g525B));
NAND2_X1 U_g8305B (.ZN(g8305B),.A2(I13285B),.A1(I13284B));
NAND2_X1 U_I5891B (.ZN(I5891B),.A2(g2057B),.A1(g750B));
NAND2_X1 U_I13273B (.ZN(I13273B),.A2(I13272B),.A1(g1918B));
NAND2_X1 U_I8480B (.ZN(I8480B),.A2(I8479B),.A1(g4455B));
NAND2_X2 U_g4144B (.ZN(g4144B),.A2(g109B),.A1(g2160B));
NAND2_X1 U_I15906B (.ZN(I15906B),.A2(g10302B),.A1(g6899B));
NAND2_X1 U_I5342B (.ZN(I5342B),.A2(I5341B),.A1(g315B));
NAND2_X1 U_I13514B (.ZN(I13514B),.A2(I13513B),.A1(g686B));
NAND2_X1 U_g8407B (.ZN(g8407B),.A2(I13523B),.A1(I13522B));
NAND2_X1 U_g4088B (.ZN(g4088B),.A2(I7225B),.A1(I7224B));
NAND2_X1 U_g4488B (.ZN(g4488B),.A2(I7877B),.A1(I7876B));
NAND2_X1 U_g7598B (.ZN(g7598B),.A2(I12138B),.A1(I12137B));
NAND3_X1 U_g3222B (.ZN(g3222B),.A3(g1834B),.A2(g1814B),.A1(g2557B));
NAND2_X1 U_I16052B (.ZN(I16052B),.A2(I16051B),.A1(g837B));
NAND2_X1 U_I12127B (.ZN(I12127B),.A2(I12126B),.A1(g6026B));
NAND2_X1 U_g10483B (.ZN(g10483B),.A2(I16088B),.A1(I16087B));
NAND2_X1 U_g8415B (.ZN(g8415B),.A2(I13561B),.A1(I13560B));
NAND2_X1 U_g11415B (.ZN(g11415B),.A2(I17290B),.A1(I17289B));
NAND2_X1 U_g6573B (.ZN(g6573B),.A2(I10509B),.A1(I10508B));
NAND2_X1 U_I5676B (.ZN(I5676B),.A2(I5675B),.A1(g1218B));
NAND2_X1 U_I6778B (.ZN(I6778B),.A2(I6777B),.A1(g2892B));
NAND2_X1 U_g9413B (.ZN(g9413B),.A2(I14614B),.A1(I14613B));
NAND2_X1 U_I8779B (.ZN(I8779B),.A2(I8778B),.A1(g4630B));
NAND2_X1 U_I5592B (.ZN(I5592B),.A2(I5591B),.A1(g1696B));
NAND4_X1 U_g8502B (.ZN(g8502B),.A4(g8366B),.A3(g591B),.A2(g605B),.A1(g2382B));
NAND2_X1 U_I15609B (.ZN(I15609B),.A2(I15607B),.A1(g10144B));
NAND2_X1 U_I15608B (.ZN(I15608B),.A2(I15607B),.A1(g10149B));
NAND3_X1 U_g3071B (.ZN(g3071B),.A3(g2382B),.A2(g2374B),.A1(g605B));
NAND2_X1 U_g10509B (.ZN(g10509B),.A2(g6023B),.A1(g10436B));
NAND2_X1 U_I17461B (.ZN(I17461B),.A2(I17459B),.A1(g11448B));
NAND2_X1 U_I13506B (.ZN(I13506B),.A2(I13504B),.A1(g8247B));
NAND2_X1 U_I5468B (.ZN(I5468B),.A2(g999B),.A1(g1245B));
NAND2_X1 U_g5219B (.ZN(g5219B),.A2(I8652B),.A1(I8651B));
NAND2_X1 U_I5677B (.ZN(I5677B),.A2(I5675B),.A1(g1223B));
NAND3_X1 U_g8826B (.ZN(g8826B),.A3(g8648B),.A2(g8737B),.A1(g8512B));
NAND2_X1 U_I17393B (.ZN(I17393B),.A2(g11414B),.A1(g11415B));
NAND2_X1 U_I5866B (.ZN(I5866B),.A2(I5865B),.A1(g2107B));
NAND2_X1 U_I12126B (.ZN(I12126B),.A2(g170B),.A1(g6026B));
NAND2_X1 U_I4978B (.ZN(I4978B),.A2(g333B),.A1(g411B));
NAND2_X1 U_g7587B (.ZN(g7587B),.A2(I12087B),.A1(I12086B));
NAND2_X1 U_g5286B (.ZN(g5286B),.A2(I8752B),.A1(I8751B));
NAND2_X1 U_g8308B (.ZN(g8308B),.A2(I13302B),.A1(I13301B));
NAND2_X1 U_I7864B (.ZN(I7864B),.A2(I7863B),.A1(g4099B));
NAND2_X1 U_I11981B (.ZN(I11981B),.A2(I11980B),.A1(g5820B));
NAND2_X1 U_I12060B (.ZN(I12060B),.A2(g1478B),.A1(g5824B));
NAND2_X1 U_g5225B (.ZN(g5225B),.A2(I8664B),.A1(I8663B));
NAND2_X1 U_g11538B (.ZN(g11538B),.A2(I17569B),.A1(I17568B));
NAND2_X1 U_I13767B (.ZN(I13767B),.A2(I13765B),.A1(g8417B));
NAND2_X1 U_g10396B (.ZN(g10396B),.A2(I15908B),.A1(I15907B));
NAND2_X1 U_I11262B (.ZN(I11262B),.A2(I11261B),.A1(g6775B));
NAND2_X1 U_I13990B (.ZN(I13990B),.A2(g8688B),.A1(g622B));
NAND2_X1 U_I6224B (.ZN(I6224B),.A2(g1346B),.A1(g2544B));
NAND2_X1 U_I5867B (.ZN(I5867B),.A2(I5865B),.A1(g2105B));
NAND2_X1 U_g2493B (.ZN(g2493B),.A2(g1840B),.A1(g1834B));
NAND2_X1 U_I5893B (.ZN(I5893B),.A2(I5891B),.A1(g2057B));
NAND3_X1 U_g3062B (.ZN(g3062B),.A3(g611B),.A2(g591B),.A1(g2369B));
NAND2_X1 U_I13521B (.ZN(I13521B),.A2(g8249B),.A1(g695B));
NAND2_X1 U_I5186B (.ZN(I5186B),.A2(I5184B),.A1(g1515B));
NAND2_X1 U_I6771B (.ZN(I6771B),.A2(I6770B),.A1(g3257B));
NAND2_X1 U_I5325B (.ZN(I5325B),.A2(I5323B),.A1(g1341B));
NAND2_X1 U_I17459B (.ZN(I17459B),.A2(g11448B),.A1(g11449B));
NAND2_X1 U_I9557B (.ZN(I9557B),.A2(g782B),.A1(g5598B));
NAND2_X1 U_g11414B (.ZN(g11414B),.A2(I17283B),.A1(I17282B));
NAND2_X1 U_I12067B (.ZN(I12067B),.A2(g139B),.A1(g6045B));
NAND2_X1 U_I12094B (.ZN(I12094B),.A2(I12092B),.A1(g1490B));
NAND2_X1 U_I4964B (.ZN(I4964B),.A2(g330B),.A1(g406B));
NAND2_X1 U_I13272B (.ZN(I13272B),.A2(g8158B),.A1(g1918B));
NAND2_X1 U_I9948B (.ZN(I9948B),.A2(I9946B),.A1(g1796B));
NAND2_X1 U_g10302B (.ZN(g10302B),.A2(I15718B),.A1(I15717B));
NAND2_X1 U_I16332B (.ZN(I16332B),.A2(I16330B),.A1(g4997B));
NAND2_X1 U_I5106B (.ZN(I5106B),.A2(I5104B),.A1(g435B));
NAND2_X1 U_g8847B (.ZN(g8847B),.A2(g8683B),.A1(g8551B));
NAND2_X1 U_g2257B (.ZN(g2257B),.A2(I5284B),.A1(I5283B));
NAND2_X1 U_I12019B (.ZN(I12019B),.A2(g166B),.A1(g6049B));
NAND2_X1 U_I15441B (.ZN(I15441B),.A2(g10007B),.A1(g10013B));
NAND2_X1 U_I11997B (.ZN(I11997B),.A2(I11995B),.A1(g127B));
NAND2_X1 U_I8739B (.ZN(I8739B),.A2(I8738B),.A1(g4607B));
NAND2_X1 U_I5461B (.ZN(I5461B),.A2(I5459B),.A1(g1003B));
NAND2_X1 U_I13766B (.ZN(I13766B),.A2(I13765B),.A1(g731B));
NAND2_X1 U_I8479B (.ZN(I8479B),.A2(g3530B),.A1(g4455B));
NAND2_X1 U_I17295B (.ZN(I17295B),.A2(g11227B),.A1(g11229B));
NAND2_X1 U_I14271B (.ZN(I14271B),.A2(I14270B),.A1(g8840B));
NAND2_X1 U_I4971B (.ZN(I4971B),.A2(g995B),.A1(g991B));
NAND2_X1 U_g8301B (.ZN(g8301B),.A2(I13267B),.A1(I13266B));
NAND2_X1 U_I6110B (.ZN(I6110B),.A2(I6109B),.A1(g2205B));
NAND2_X1 U_g10482B (.ZN(g10482B),.A2(I16081B),.A1(I16080B));
NAND2_X1 U_g10779B (.ZN(g10779B),.A2(I16469B),.A1(I16468B));
NAND2_X1 U_I6762B (.ZN(I6762B),.A2(I6760B),.A1(g1448B));
NAND2_X1 U_I17289B (.ZN(I17289B),.A2(I17288B),.A1(g11225B));
NAND2_X1 U_I5315B (.ZN(I5315B),.A2(g1027B),.A1(g1032B));
NAND2_X1 U_I17288B (.ZN(I17288B),.A2(g11223B),.A1(g11225B));
NAND2_X1 U_I13859B (.ZN(I13859B),.A2(I13857B),.A1(g1448B));
NAND2_X1 U_g7548B (.ZN(g7548B),.A2(I11982B),.A1(I11981B));
NAND2_X1 U_I13858B (.ZN(I13858B),.A2(I13857B),.A1(g8270B));
NAND2_X1 U_I11996B (.ZN(I11996B),.A2(I11995B),.A1(g6035B));
NAND3_X1 U_g8743B (.ZN(g8743B),.A3(I9265B),.A2(I9273B),.A1(g8617B));
NAND2_X1 U_I5880B (.ZN(I5880B),.A2(I5878B),.A1(g2115B));
NAND2_X1 U_g10513B (.ZN(g10513B),.A2(g5345B),.A1(g10441B));
NAND2_X1 U_g8411B (.ZN(g8411B),.A2(I13539B),.A1(I13538B));
NAND2_X1 U_I8626B (.ZN(I8626B),.A2(I8624B),.A1(g511B));
NAND2_X1 U_g10505B (.ZN(g10505B),.A2(g5938B),.A1(g10432B));
NAND2_X1 U_I5612B (.ZN(I5612B),.A2(I5611B),.A1(g1280B));
NAND2_X1 U_g4821B (.ZN(g4821B),.A2(I8180B),.A1(I8179B));
NAND2_X1 U_I12076B (.ZN(I12076B),.A2(I12074B),.A1(g174B));
NAND2_X1 U_I12085B (.ZN(I12085B),.A2(g1470B),.A1(g5842B));
NAND2_X1 U_g7567B (.ZN(g7567B),.A2(I12021B),.A1(I12020B));
NAND2_X1 U_I5128B (.ZN(I5128B),.A2(I5126B),.A1(g1389B));
NAND2_X1 U_I6489B (.ZN(I6489B),.A2(I6487B),.A1(g1227B));
NAND2_X1 U_g7593B (.ZN(g7593B),.A2(I12115B),.A1(I12114B));
NAND2_X1 U_I8778B (.ZN(I8778B),.A2(g1137B),.A1(g4630B));
NAND2_X1 U_g10149B (.ZN(g10149B),.A2(I15443B),.A1(I15442B));
NAND2_X1 U_I13902B (.ZN(I13902B),.A2(I13900B),.A1(g1428B));
NAND2_X1 U_I13301B (.ZN(I13301B),.A2(I13300B),.A1(g1936B));
NAND2_X1 U_g3215B (.ZN(g3215B),.A2(g1822B),.A1(g2564B));
NAND4_X1 U_g7996B (.ZN(g7996B),.A4(FE_OFN96_g2169B),.A3(g7562B),.A2(g7574B),.A1(FE_OFN88_g2178B));
NAND2_X1 U_I4985B (.ZN(I4985B),.A2(g1003B),.A1(g999B));
NAND2_X1 U_I14444B (.ZN(I14444B),.A2(I14442B),.A1(g1834B));
NAND4_X1 U_g8000B (.ZN(g8000B),.A4(g7550B),.A3(g7562B),.A2(g7574B),.A1(FE_OFN88_g2178B));
NAND2_X1 U_I5166B (.ZN(I5166B),.A2(I5164B),.A1(g1499B));
NAND2_X1 U_I17460B (.ZN(I17460B),.A2(I17459B),.A1(g11449B));
NAND2_X1 U_g3008B (.ZN(g3008B),.A2(g878B),.A1(g2444B));
NAND2_X1 U_I6836B (.ZN(I6836B),.A2(g806B),.A1(g3287B));
NAND2_X1 U_I5529B (.ZN(I5529B),.A2(I5528B),.A1(g1265B));
NAND2_X1 U_g10229B (.ZN(g10229B),.A2(I15609B),.A1(I15608B));
NAND2_X1 U_I13661B (.ZN(I13661B),.A2(I13659B),.A1(g8322B));
NAND2_X1 U_I13895B (.ZN(I13895B),.A2(I13893B),.A1(g1436B));
NAND2_X1 U_g2303B (.ZN(g2303B),.A2(I5343B),.A1(I5342B));
NAND2_X1 U_I12039B (.ZN(I12039B),.A2(I12038B),.A1(g5847B));
NAND2_X1 U_g5592B (.ZN(g5592B),.A2(I9008B),.A1(I9007B));
NAND2_X1 U_I12038B (.ZN(I12038B),.A2(g1466B),.A1(g5847B));
NAND2_X1 U_g3322B (.ZN(g3322B),.A2(I6489B),.A1(I6488B));
NAND2_X1 U_I8561B (.ZN(I8561B),.A2(g491B),.A1(g4227B));
NAND2_X1 U_I8527B (.ZN(I8527B),.A2(g481B),.A1(g4879B));
NAND2_X1 U_I12143B (.ZN(I12143B),.A2(g158B),.A1(g6000B));
NAND2_X1 U_I5619B (.ZN(I5619B),.A2(I5618B),.A1(g1766B));
NAND2_X1 U_g10386B (.ZN(g10386B),.A2(I15880B),.A1(I15879B));
NAND2_X1 U_I11980B (.ZN(I11980B),.A2(g1482B),.A1(g5820B));
NAND2_X1 U_I6837B (.ZN(I6837B),.A2(I6836B),.A1(g3287B));
NAND2_X1 U_I4973B (.ZN(I4973B),.A2(I4971B),.A1(g995B));
NAND2_X1 U_I13888B (.ZN(I13888B),.A2(I13886B),.A1(g1440B));
NAND2_X1 U_g7558B (.ZN(g7558B),.A2(I12004B),.A1(I12003B));
NAND2_X1 U_I17494B (.ZN(I17494B),.A2(I17492B),.A1(g3623B));
NAND2_X1 U_g11491B (.ZN(g11491B),.A2(I17494B),.A1(I17493B));
NAND2_X1 U_I16045B (.ZN(I16045B),.A2(I16044B),.A1(g833B));
NAND2_X1 U_I7684B (.ZN(I7684B),.A2(I7683B),.A1(g1023B));
NAND2_X1 U_g4130B (.ZN(g4130B),.A2(g2518B),.A1(FE_OFN352_g109B));
NAND2_X1 U_I8771B (.ZN(I8771B),.A2(I8770B),.A1(g4619B));
NAND2_X1 U_I13546B (.ZN(I13546B),.A2(I13544B),.A1(g8259B));
NAND2_X1 U_I13089B (.ZN(I13089B),.A2(g1840B),.A1(g8006B));
NAND2_X1 U_g2117B (.ZN(g2117B),.A2(I5025B),.A1(I5024B));
NAND2_X1 U_g5119B (.ZN(g5119B),.A2(I8515B),.A1(I8514B));
NAND2_X1 U_g5319B (.ZN(g5319B),.A2(I8805B),.A1(I8804B));
NAND2_X1 U_I15899B (.ZN(I15899B),.A2(I15898B),.A1(g857B));
NAND2_X1 U_I5606B (.ZN(I5606B),.A2(I5604B),.A1(g1153B));
NAND2_X1 U_I15898B (.ZN(I15898B),.A2(g10359B),.A1(g857B));
NAND2_X1 U_I16032B (.ZN(I16032B),.A2(I16030B),.A1(g10430B));
NAND2_X1 U_I17401B (.ZN(I17401B),.A2(I17400B),.A1(g11418B));
NAND2_X1 U_I13659B (.ZN(I13659B),.A2(g8322B),.A1(g1945B));
NAND2_X1 U_I8738B (.ZN(I8738B),.A2(g1121B),.A1(g4607B));
NAND2_X1 U_I13250B (.ZN(I13250B),.A2(I13248B),.A1(g8148B));
NAND2_X1 U_I15718B (.ZN(I15718B),.A2(I15716B),.A1(g10229B));
NAND2_X1 U_I9008B (.ZN(I9008B),.A2(I9006B),.A1(FE_OFN252_g1791B));
NAND2_X1 U_I6176B (.ZN(I6176B),.A2(g197B),.A1(g2177B));
NAND2_X1 U_I7865B (.ZN(I7865B),.A2(I7863B),.A1(g774B));
NAND2_X1 U_g5274B (.ZN(g5274B),.A2(I8730B),.A1(I8729B));
NAND2_X1 U_I5341B (.ZN(I5341B),.A2(g426B),.A1(g315B));
NAND2_X1 U_I17305B (.ZN(I17305B),.A2(g11231B),.A1(g11232B));
NAND2_X1 U_I17053B (.ZN(I17053B),.A2(I17051B),.A1(g11249B));
NAND2_X1 U_g5125B (.ZN(g5125B),.A2(I8529B),.A1(I8528B));
NAND2_X1 U_I12216B (.ZN(I12216B),.A2(I12214B),.A1(g2518B));
NAND2_X1 U_I6225B (.ZN(I6225B),.A2(I6224B),.A1(g2544B));
NAND2_X1 U_I5879B (.ZN(I5879B),.A2(I5878B),.A1(g2120B));
NAND2_X1 U_g3221B (.ZN(g3221B),.A2(g2564B),.A1(g1834B));
NAND2_X1 U_I14270B (.ZN(I14270B),.A2(g1822B),.A1(g8840B));
NAND2_X1 U_I6124B (.ZN(I6124B),.A2(g1419B),.A1(g2215B));
NAND2_X1 U_I6324B (.ZN(I6324B),.A2(I6322B),.A1(g1864B));
NAND2_X1 U_I13867B (.ZN(I13867B),.A2(g1403B),.A1(g8264B));
NAND2_X1 U_I13894B (.ZN(I13894B),.A2(I13893B),.A1(g8266B));
NAND2_X1 U_I6469B (.ZN(I6469B),.A2(I6467B),.A1(g2479B));
NAND2_X1 U_I8663B (.ZN(I8663B),.A2(I8662B),.A1(g4286B));
NAND2_X1 U_g7523B (.ZN(g7523B),.A2(I11909B),.A1(I11908B));
NAND2_X1 U_I6177B (.ZN(I6177B),.A2(I6176B),.A1(g2177B));
NAND2_X1 U_g5187B (.ZN(g5187B),.A2(I8591B),.A1(I8590B));
NAND2_X1 U_I6287B (.ZN(I6287B),.A2(g981B),.A1(g2091B));
NAND2_X1 U_I8762B (.ZN(I8762B),.A2(I8761B),.A1(g4616B));
NAND2_X1 U_I15871B (.ZN(I15871B),.A2(I15870B),.A1(g10291B));
NAND3_X1 U_g8840B (.ZN(g8840B),.A3(g8551B),.A2(g8541B),.A1(g8542B));
NAND2_X1 U_g2250B (.ZN(g2250B),.A2(I5265B),.A1(I5264B));
NAND2_X1 U_I8590B (.ZN(I8590B),.A2(I8589B),.A1(g4251B));
NAND2_X1 U_I6199B (.ZN(I6199B),.A2(g766B),.A1(g2525B));
NAND2_X1 U_I14218B (.ZN(I14218B),.A2(I14216B),.A1(g605B));
NAND2_X1 U_g8190B (.ZN(g8190B),.A2(g7978B),.A1(g6027B));
NAND2_X1 U_I5284B (.ZN(I5284B),.A2(I5282B),.A1(g762B));
NAND2_X1 U_I17485B (.ZN(I17485B),.A2(g11474B),.A1(g11233B));
NAND2_X1 U_I4965B (.ZN(I4965B),.A2(I4964B),.A1(g406B));
NAND2_X1 U_I5591B (.ZN(I5591B),.A2(g1703B),.A1(g1696B));
NAND2_X1 U_g8501B (.ZN(g8501B),.A2(g8366B),.A1(g3760B));
NAND2_X1 U_I15451B (.ZN(I15451B),.A2(g10019B),.A1(g10025B));
NAND2_X1 U_g8942B (.ZN(g8942B),.A2(FE_OFN200_g4921B),.A1(g8823B));
NAND2_X1 U_I13877B (.ZN(I13877B),.A2(I13876B),.A1(g8269B));
NAND2_X1 U_g7269B (.ZN(g7269B),.A2(I11510B),.A1(I11509B));
NAND2_X1 U_I4996B (.ZN(I4996B),.A2(I4995B),.A1(g416B));
NAND2_X1 U_I6144B (.ZN(I6144B),.A2(I6143B),.A1(g1976B));
NAND2_X1 U_I17567B (.ZN(I17567B),.A2(g1610B),.A1(g11496B));
NAND2_X1 U_g7572B (.ZN(g7572B),.A2(I12040B),.A1(I12039B));
NAND2_X1 U_I6207B (.ZN(I6207B),.A2(g802B),.A1(g5188B));
NAND2_X1 U_I14277B (.ZN(I14277B),.A2(g1828B),.A1(g8847B));
NAND2_X1 U_I16059B (.ZN(I16059B),.A2(I16058B),.A1(g841B));
NAND2_X1 U_I16025B (.ZN(I16025B),.A2(I16023B),.A1(FE_OFN253_g1786B));
NAND2_X1 U_I8563B (.ZN(I8563B),.A2(I8561B),.A1(g491B));
NAND2_X1 U_g3524B (.ZN(g3524B),.A2(g3221B),.A1(g3209B));
NAND2_X1 U_I16058B (.ZN(I16058B),.A2(g10441B),.A1(g841B));
NAND2_X1 U_I5204B (.ZN(I5204B),.A2(I5202B),.A1(g374B));
NAND2_X1 U_I6488B (.ZN(I6488B),.A2(I6487B),.A1(g2306B));
NAND4_X1 U_g3818B (.ZN(g3818B),.A4(g3003B),.A3(g2310B),.A2(g3071B),.A1(g3056B));
NAND2_X1 U_I16044B (.ZN(I16044B),.A2(g10432B),.A1(g833B));
NAND2_X1 U_g3717B (.ZN(g3717B),.A2(I6881B),.A1(I6880B));
NAND2_X1 U_I13077B (.ZN(I13077B),.A2(I13076B),.A1(g1872B));
NAND2_X1 U_g10043B (.ZN(g10043B),.A2(I15258B),.A1(I15257B));
NAND2_X1 U_I11280B (.ZN(I11280B),.A2(I11278B),.A1(g6485B));
NAND2_X1 U_I6825B (.ZN(I6825B),.A2(g770B),.A1(g3281B));
NAND2_X1 U_I4997B (.ZN(I4997B),.A2(I4995B),.A1(g309B));
NAND2_X1 U_I13300B (.ZN(I13300B),.A2(g8162B),.A1(g1936B));
NAND2_X1 U_I5323B (.ZN(I5323B),.A2(g1341B),.A1(g1336B));
NAND2_X1 U_I6136B (.ZN(I6136B),.A2(g378B),.A1(g2496B));
NAND2_X1 U_g5935B (.ZN(g5935B),.A2(I9559B),.A1(I9558B));
NAND2_X1 U_I5528B (.ZN(I5528B),.A2(g1015B),.A1(g1265B));
NAND2_X1 U_I6806B (.ZN(I6806B),.A2(I6805B),.A1(g3268B));
NAND2_X1 U_I5530B (.ZN(I5530B),.A2(I5528B),.A1(g1015B));
NAND2_X1 U_g10886B (.ZN(g10886B),.A2(g10805B),.A1(g10807B));
NAND2_X1 U_g3106B (.ZN(g3106B),.A2(I6324B),.A1(I6323B));
NAND2_X1 U_I13876B (.ZN(I13876B),.A2(g1444B),.A1(g8269B));
NAND2_X1 U_I6322B (.ZN(I6322B),.A2(g1864B),.A1(g2050B));
NAND2_X1 U_g3061B (.ZN(g3061B),.A2(g2374B),.A1(g611B));
NAND2_X1 U_g2439B (.ZN(g2439B),.A2(g1828B),.A1(g1814B));
NAND4_X1 U_g7947B (.ZN(g7947B),.A4(g7550B),.A3(FE_OFN91_g2172B),.A2(g7574B),.A1(g6941B));
NAND2_X1 U_I9576B (.ZN(I9576B),.A2(I9574B),.A1(g818B));
NAND2_X1 U_I13660B (.ZN(I13660B),.A2(I13659B),.A1(g1945B));
NAND2_X1 U_g3200B (.ZN(g3200B),.A2(g2061B),.A1(g1822B));
NAND2_X1 U_g4374B (.ZN(g4374B),.A2(I7685B),.A1(I7684B));
NAND2_X1 U_I11916B (.ZN(I11916B),.A2(I11914B),.A1(g1494B));
NAND2_X1 U_I5372B (.ZN(I5372B),.A2(I5371B),.A1(g971B));
NAND2_X1 U_g3003B (.ZN(g3003B),.A2(g2399B),.A1(g599B));
NAND2_X1 U_g8627B (.ZN(g8627B),.A2(I13888B),.A1(I13887B));
NAND2_X1 U_I5618B (.ZN(I5618B),.A2(FE_OFN247_g1771B),.A1(g1766B));
NAND2_X1 U_I6137B (.ZN(I6137B),.A2(I6136B),.A1(g2496B));
NAND2_X1 U_I5343B (.ZN(I5343B),.A2(I5341B),.A1(g426B));
NAND2_X1 U_I5282B (.ZN(I5282B),.A2(g762B),.A1(g758B));
NAND2_X1 U_I13307B (.ZN(I13307B),.A2(g617B),.A1(g8190B));
NAND2_X1 U_I13076B (.ZN(I13076B),.A2(g7963B),.A1(g1872B));
NAND2_X1 U_I6807B (.ZN(I6807B),.A2(I6805B),.A1(g471B));
NAND2_X1 U_I11243B (.ZN(I11243B),.A2(I11241B),.A1(g790B));
NAND2_X1 U_I17585B (.ZN(I17585B),.A2(I17584B),.A1(g11217B));
NAND2_X1 U_I12137B (.ZN(I12137B),.A2(I12136B),.A1(g6038B));
NAND2_X1 U_I7564B (.ZN(I7564B),.A2(I7562B),.A1(g654B));
NAND2_X1 U_g2970B (.ZN(g2970B),.A2(I6201B),.A1(I6200B));
NAND2_X1 U_g10144B (.ZN(g10144B),.A2(I15432B),.A1(I15431B));
NAND2_X1 U_I8788B (.ZN(I8788B),.A2(I8786B),.A1(g1141B));
NAND2_X1 U_g7054B (.ZN(g7054B),.A2(I11243B),.A1(I11242B));
NAND2_X1 U_I17052B (.ZN(I17052B),.A2(I17051B),.A1(g10923B));
NAND2_X1 U_g2120B (.ZN(g2120B),.A2(I5036B),.A1(I5035B));
NAND2_X1 U_g8616B (.ZN(g8616B),.A2(I13869B),.A1(I13868B));
NAND2_X1 U_I5202B (.ZN(I5202B),.A2(g374B),.A1(g369B));
NAND2_X1 U_I16088B (.ZN(I16088B),.A2(I16086B),.A1(g10430B));
NAND2_X1 U_I16024B (.ZN(I16024B),.A2(I16023B),.A1(g10438B));
NAND2_X1 U_g11490B (.ZN(g11490B),.A2(I17487B),.A1(I17486B));
NAND2_X1 U_I5518B (.ZN(I5518B),.A2(I5516B),.A1(g1019B));
NAND3_X1 U_g5118B (.ZN(g5118B),.A3(g4073B),.A2(g4806B),.A1(g2439B));
NAND2_X1 U_I12021B (.ZN(I12021B),.A2(I12019B),.A1(g166B));
NOR2_X1 U_g6392B (.ZN(g6392B),.A2(g5938B),.A1(g5859B));
NOR2_X1 U_g5938B (.ZN(g5938B),.A2(FE_OFN349_I6424B),.A1(g2273B));
NOR2_X1 U_g2478B (.ZN(g2478B),.A2(g1737B),.A1(g1610B));
NOR4_X1 U_g4278B (.ZN(g4278B),.A4(g3776B),.A3(FE_OFN254_g461B),.A2(FE_OFN248_g466B),.A1(g3800B));
NOR2_X1 U_g10383B (.ZN(g10383B),.A2(g3348B),.A1(I15514B));
NOR2_X1 U_g3118B (.ZN(g3118B),.A2(g2514B),.A1(g2521B));
NOR2_X1 U_g9815B (.ZN(g9815B),.A2(FE_OFN67_g9367B),.A1(FE_OFN68_g9392B));
NOR2_X1 U_g11077B (.ZN(g11077B),.A2(g10971B),.A1(g10970B));
NOR3_X1 U_g3879B (.ZN(g3879B),.A3(g2353B),.A2(g2354B),.A1(g3141B));
NOR2_X1 U_g10285B (.ZN(g10285B),.A2(FE_OFN350_g3121B),.A1(I15287B));
NOR2_X1 U_g11480B (.ZN(g11480B),.A2(g4567B),.A1(g11456B));
NOR2_X1 U_g4076B (.ZN(g4076B),.A2(I5254B),.A1(g1707B));
NOR2_X1 U_g10570B (.ZN(g10570B),.A2(g10324B),.A1(g10485B));
NOR2_X1 U_g10239B (.ZN(g10239B),.A2(I15287B),.A1(g9317B));
NOR2_X1 U_g10594B (.ZN(g10594B),.A2(g10521B),.A1(g10480B));
NOR2_X1 U_g9426B (.ZN(g9426B),.A2(FE_OFN50_g9030B),.A1(FE_OFN54_g9052B));
NOR2_X1 U_g10382B (.ZN(g10382B),.A2(g3348B),.A1(I15507B));
NOR4_X1 U_g4672B (.ZN(g4672B),.A4(g3479B),.A3(g1104B),.A2(g1107B),.A1(g3501B));
NOR2_X1 U_g5360B (.ZN(g5360B),.A2(FE_OFN308_I6424B),.A1(g105B));
NOR4_X1 U_g9387B (.ZN(g9387B),.A4(I14779B),.A3(g9223B),.A2(g9240B),.A1(g9010B));
NOR2_X1 U_g10438B (.ZN(g10438B),.A2(FE_OFN160_I6424B),.A1(I15500B));
NOR4_X1 U_g4613B (.ZN(g4613B),.A4(g1101B),.A3(g1104B),.A2(g3491B),.A1(FE_OFN240_g1110B));
NOR4_X1 U_g9391B (.ZN(g9391B),.A4(I14602B),.A3(FE_OFN39_g9223B),.A2(FE_OFN40_g9240B),.A1(g9010B));
NOR3_X1 U_g4572B (.ZN(g4572B),.A3(g3628B),.A2(g3408B),.A1(g3419B));
NOR3_X1 U_g9757B (.ZN(g9757B),.A3(FE_OFN72_g9292B),.A2(FE_OFN62_g9274B),.A1(FE_OFN32_g9454B));
NOR4_X1 U_g9874B (.ZN(g9874B),.A4(I15033B),.A3(g9579B),.A2(FE_OFN64_g9536B),.A1(g9519B));
NOR2_X1 U_g9654B (.ZN(g9654B),.A2(FE_OFN53_g9173B),.A1(FE_OFN46_g9125B));
NOR4_X1 U_g9880B (.ZN(g9880B),.A4(I15051B),.A3(g9579B),.A2(FE_OFN64_g9536B),.A1(g9751B));
NOR4_X1 U_g4873B (.ZN(g4873B),.A4(g3776B),.A3(FE_OFN254_g461B),.A2(FE_OFN248_g466B),.A1(FE_OFN250_g471B));
NOR2_X1 U_g2807B (.ZN(g2807B),.A2(g3629B),.A1(FE_OFN266_g18B));
NOR2_X1 U_g10441B (.ZN(g10441B),.A2(FE_OFN160_I6424B),.A1(I15510B));
NOR4_X1 U_g4639B (.ZN(g4639B),.A4(g1101B),.A3(g1104B),.A2(g1107B),.A1(g3501B));
NOR2_X1 U_g10435B (.ZN(g10435B),.A2(g3744B),.A1(I15510B));
NOR2_X1 U_g10849B (.ZN(g10849B),.A2(g2459B),.A1(g10739B));
NOR4_X1 U_g9606B (.ZN(g9606B),.A4(FE_OFN48_g9151B),.A3(FE_OFN52_g9173B),.A2(FE_OFN51_g9111B),.A1(FE_OFN45_g9125B));
NOR4_X1 U_g9879B (.ZN(g9879B),.A4(I15048B),.A3(g9563B),.A2(FE_OFN64_g9536B),.A1(g9747B));
NOR2_X1 U_g9506B (.ZN(g9506B),.A2(FE_OFN49_g9030B),.A1(FE_OFN56_g9052B));
NOR2_X1 U_g6155B (.ZN(g6155B),.A2(I5254B),.A1(g4974B));
NOR2_X1 U_g6355B (.ZN(g6355B),.A2(g6023B),.A1(g6032B));
NOR2_X1 U_g9591B (.ZN(g9591B),.A2(FE_OFN47_g9151B),.A1(FE_OFN44_g9125B));
NOR2_X1 U_g10359B (.ZN(g10359B),.A2(FE_OFN308_I6424B),.A1(I15290B));
NOR2_X1 U_g10434B (.ZN(g10434B),.A2(FE_OFN349_I6424B),.A1(I15514B));
NOR2_X1 U_g10291B (.ZN(g10291B),.A2(FE_OFN308_I6424B),.A1(I15287B));
NOR4_X1 U_g4227B (.ZN(g4227B),.A4(g2579B),.A3(FE_OFN254_g461B),.A2(g3793B),.A1(FE_OFN250_g471B));
NOR4_X1 U_g9667B (.ZN(g9667B),.A4(FE_OFN47_g9151B),.A3(FE_OFN52_g9173B),.A2(FE_OFN51_g9111B),.A1(FE_OFN45_g9125B));
NOR2_X1 U_g10563B (.ZN(g10563B),.A2(g10322B),.A1(g10484B));
NOR2_X1 U_g10324B (.ZN(g10324B),.A2(I15365B),.A1(g9317B));
NOR3_X1 U_g4455B (.ZN(g4455B),.A3(g3408B),.A2(g3419B),.A1(g3543B));
NOR4_X1 U_g9878B (.ZN(g9878B),.A4(I15045B),.A3(g9579B),.A2(FE_OFN64_g9536B),.A1(g9754B));
NOR2_X1 U_g10360B (.ZN(g10360B),.A2(FE_OFN350_g3121B),.A1(I15290B));
NOR4_X1 U_g9882B (.ZN(g9882B),.A4(I15057B),.A3(g9563B),.A2(FE_OFN64_g9536B),.A1(g9747B));
NOR4_X1 U_g4605B (.ZN(g4605B),.A4(g1101B),.A3(g3485B),.A2(g1107B),.A1(FE_OFN240_g1110B));
NOR2_X1 U_g10562B (.ZN(g10562B),.A2(g10529B),.A1(g10483B));
NOR2_X1 U_g5780B (.ZN(g5780B),.A2(FE_OFN200_g4921B),.A1(g3092B));
NOR2_X1 U_g10385B (.ZN(g10385B),.A2(g3348B),.A1(I15510B));
NOR4_X1 U_g4601B (.ZN(g4601B),.A4(g3479B),.A3(g1104B),.A2(g1107B),.A1(FE_OFN240_g1110B));
NOR2_X1 U_g5573B (.ZN(g5573B),.A2(g4432B),.A1(g4117B));
NOR2_X1 U_g5999B (.ZN(g5999B),.A2(FE_OFN349_I6424B),.A1(g2271B));
NOR3_X1 U_g9759B (.ZN(g9759B),.A3(FE_OFN71_g9292B),.A2(g9274B),.A1(g9454B));
NOR2_X1 U_g6037B (.ZN(g6037B),.A2(FE_OFN350_g3121B),.A1(g2297B));
NOR2_X1 U_g5034B (.ZN(g5034B),.A2(g3967B),.A1(g3524B));
NOR4_X1 U_g9881B (.ZN(g9881B),.A4(I15054B),.A3(g9579B),.A2(FE_OFN64_g9536B),.A1(g9516B));
NOR3_X1 U_g4276B (.ZN(g4276B),.A3(g2500B),.A2(g3261B),.A1(g4065B));
NOR4_X1 U_g4616B (.ZN(g4616B),.A4(g3479B),.A3(g1104B),.A2(g3491B),.A1(FE_OFN240_g1110B));
NOR2_X1 U_g10363B (.ZN(g10363B),.A2(FE_OFN308_I6424B),.A1(I15365B));
NOR2_X1 U_g2862B (.ZN(g2862B),.A2(g2305B),.A1(g2315B));
NOR3_X1 U_g9758B (.ZN(g9758B),.A3(FE_OFN71_g9292B),.A2(FE_OFN62_g9274B),.A1(FE_OFN32_g9454B));
NOR3_X1 U_g9589B (.ZN(g9589B),.A3(FE_OFN48_g9151B),.A2(FE_OFN52_g9173B),.A1(FE_OFN45_g9125B));
NOR2_X1 U_g9803B (.ZN(g9803B),.A2(g9367B),.A1(FE_OFN69_g9392B));
NOR2_X1 U_g10430B (.ZN(g10430B),.A2(FE_OFN349_I6424B),.A1(I15503B));
NOR2_X1 U_g10362B (.ZN(g10362B),.A2(g3744B),.A1(I15290B));
NOR2_X1 U_g2791B (.ZN(g2791B),.A2(g750B),.A1(g2187B));
NOR4_X1 U_g9605B (.ZN(g9605B),.A4(FE_OFN48_g9151B),.A3(FE_OFN52_g9173B),.A2(FE_OFN51_g9111B),.A1(FE_OFN46_g9125B));
NOR2_X1 U_g10436B (.ZN(g10436B),.A2(FE_OFN349_I6424B),.A1(I15510B));
NOR4_X1 U_g5556B (.ZN(g5556B),.A4(g2031B),.A3(g2299B),.A2(FE_OFN238_g1781B),.A1(g4787B));
NOR4_X1 U_g4286B (.ZN(g4286B),.A4(g2579B),.A3(g3784B),.A2(FE_OFN248_g466B),.A1(g3800B));
NOR2_X1 U_g4974B (.ZN(g4974B),.A2(g3714B),.A1(g4502B));
NOR2_X1 U_g9423B (.ZN(g9423B),.A2(FE_OFN49_g9030B),.A1(FE_OFN54_g9052B));
NOR2_X1 U_g5350B (.ZN(g5350B),.A2(FE_OFN160_I6424B),.A1(g3070B));
NOR4_X1 U_g2459B (.ZN(g2459B),.A4(g1648B),.A3(g1651B),.A2(g1642B),.A1(g1645B));
NOR2_X1 U_g10381B (.ZN(g10381B),.A2(g3348B),.A1(I15503B));
NOR4_X1 U_g4259B (.ZN(g4259B),.A4(g3776B),.A3(g3784B),.A2(g3793B),.A1(FE_OFN250_g471B));
NOR2_X1 U_g10522B (.ZN(g10522B),.A2(g10239B),.A1(g10401B));
NOR2_X1 U_g5392B (.ZN(g5392B),.A2(FE_OFN160_I6424B),.A1(g3086B));
NOR3_X1 U_g4122B (.ZN(g4122B),.A3(g2538B),.A2(g2410B),.A1(g3291B));
NOR2_X1 U_g6023B (.ZN(g6023B),.A2(FE_OFN160_I6424B),.A1(g2275B));
NOR2_X1 U_g3462B (.ZN(g3462B),.A2(g2795B),.A1(g2187B));
NOR4_X1 U_g4218B (.ZN(g4218B),.A4(g3776B),.A3(g3784B),.A2(FE_OFN248_g466B),.A1(FE_OFN250_g471B));
NOR4_X1 U_g4267B (.ZN(g4267B),.A4(g2579B),.A3(FE_OFN254_g461B),.A2(FE_OFN248_g466B),.A1(g3800B));
NOR4_X1 U_g4677B (.ZN(g4677B),.A4(g1101B),.A3(g3485B),.A2(g1107B),.A1(g3501B));
NOR2_X1 U_g9646B (.ZN(g9646B),.A2(FE_OFN47_g9151B),.A1(FE_OFN45_g9125B));
NOR2_X1 U_g2863B (.ZN(g2863B),.A2(g2309B),.A1(g2316B));
NOR2_X1 U_g6032B (.ZN(g6032B),.A2(FE_OFN349_I6424B),.A1(g3008B));
NOR4_X1 U_g9647B (.ZN(g9647B),.A4(FE_OFN48_g9151B),.A3(FE_OFN53_g9173B),.A2(FE_OFN51_g9111B),.A1(FE_OFN46_g9125B));
NOR2_X1 U_g5859B (.ZN(g5859B),.A2(FE_OFN349_I6424B),.A1(g2987B));
NOR2_X1 U_g10433B (.ZN(g10433B),.A2(g3744B),.A1(I15514B));
NOR4_X1 U_g4251B (.ZN(g4251B),.A4(g2579B),.A3(g3784B),.A2(g3793B),.A1(FE_OFN250_g471B));
NOR4_X1 U_g9876B (.ZN(g9876B),.A4(I15054B),.A3(FE_OFN56_g9052B),.A2(FE_OFN280_g9536B),.A1(g9522B));
NOR2_X1 U_g8303B (.ZN(g8303B),.A2(g4811B),.A1(g8209B));
NOR2_X1 U_g10429B (.ZN(g10429B),.A2(g3744B),.A1(I15503B));
NOR2_X1 U_g10428B (.ZN(g10428B),.A2(g3121B),.A1(I15503B));
NOR4_X1 U_g4234B (.ZN(g4234B),.A4(g3776B),.A3(FE_OFN254_g461B),.A2(g3793B),.A1(FE_OFN250_g471B));
NOR4_X1 U_g9877B (.ZN(g9877B),.A4(I15048B),.A3(g9569B),.A2(FE_OFN64_g9536B),.A1(g9512B));
NOR2_X1 U_g5186B (.ZN(g5186B),.A2(FE_OFN223_g4401B),.A1(g2047B));
NOR4_X1 U_g4619B (.ZN(g4619B),.A4(g1101B),.A3(g3485B),.A2(g3491B),.A1(FE_OFN240_g1110B));
NOR2_X1 U_g10432B (.ZN(g10432B),.A2(FE_OFN349_I6424B),.A1(I15507B));
NOR2_X1 U_g5345B (.ZN(g5345B),.A2(FE_OFN350_g3121B),.A1(g2067B));
NOR2_X1 U_g5763B (.ZN(g5763B),.A2(g5345B),.A1(g5350B));
NOR4_X1 U_g4879B (.ZN(g4879B),.A4(g2579B),.A3(g3784B),.A2(FE_OFN248_g466B),.A1(FE_OFN250_g471B));
NOR4_X1 U_g4607B (.ZN(g4607B),.A4(g3479B),.A3(g3485B),.A2(g1107B),.A1(FE_OFN240_g1110B));
NOR2_X1 U_g3107B (.ZN(g3107B),.A2(g2499B),.A1(g2501B));
NOR2_X1 U_g10322B (.ZN(g10322B),.A2(I15500B),.A1(g9317B));
NOR4_X1 U_g4630B (.ZN(g4630B),.A4(g3479B),.A3(g3485B),.A2(g3491B),.A1(FE_OFN240_g1110B));
NOR2_X1 U_g10364B (.ZN(g10364B),.A2(g3744B),.A1(I15507B));
SDFF_X1 U_g1289B (.Q(g1289B),.SE(test_seB),.SI(test_siB),.D(g4556B),.CK(CKB));
SDFF_X1 U_g1882B (.Q(g1882B),.SE(test_seB),.SI(g1289B),.D(g8943B),.CK(CKB));
SDFF_X1 U_g312B (.Q(g312B),.SE(test_seB),.SI(g1882B),.D(g255B),.CK(CKB));
SDFF_X1 U_g452B (.Q(g452B),.SE(test_seB),.SI(g312B),.D(g11257B),.CK(CKB));
SDFF_X1 U_g123B (.Q(g123B),.SE(test_seB),.SI(g452B),.D(g7032B),.CK(CKB));
SDFF_X1 U_g207B (.Q(g207B),.SE(test_seB),.SI(g123B),.D(g6830B),.CK(CKB));
SDFF_X1 U_g713B (.Q(g713B),.SE(test_seB),.SI(g207B),.D(g8920B),.CK(CKB));
SDFF_X1 U_g1153B (.Q(g1153B),.SE(test_seB),.SI(g713B),.D(g4340B),.CK(CKB));
SDFF_X1 U_g1209B (.Q(g1209B),.SE(test_seB),.SI(g1153B),.D(g10732B),.CK(CKB));
SDFF_X1 U_g1744B (.Q(g1744B),.SE(test_seB),.SI(g1209B),.D(g4239B),.CK(CKB));
SDFF_X1 U_g1558B (.Q(g1558B),.SE(test_seB),.SI(g1744B),.D(g6538B),.CK(CKB));
SDFF_X1 U_g695B (.Q(g695B),.SE(test_seB),.SI(g1558B),.D(g8887B),.CK(CKB));
SDFF_X1 U_g461B (.Q(g461B),.SE(test_seB),.SI(g695B),.D(g11372B),.CK(CKB));
SDFF_X1 U_g940B (.Q(g940B),.SE(test_seB),.SI(g461B),.D(g8260B),.CK(CKB));
SDFF_X1 U_g976B (.Q(g976B),.SE(test_seB),.SI(g940B),.D(g11391B),.CK(CKB));
SDFF_X1 U_g709B (.Q(g709B),.SE(test_seB),.SI(g976B),.D(g8432B),.CK(CKB));
SDFF_X1 U_g1092B (.Q(g1092B),.SE(test_seB),.SI(g709B),.D(g6088B),.CK(CKB));
SDFF_X1 U_g1574B (.Q(g1574B),.SE(test_seB),.SI(g1092B),.D(g6478B),.CK(CKB));
SDFF_X1 U_g1864B (.Q(g1864B),.SE(test_seB),.SI(g1574B),.D(g6795B),.CK(CKB));
SDFF_X1 U_g369B (.Q(g369B),.SE(test_seB),.SI(g1864B),.D(g11320B),.CK(CKB));
SDFF_X1 U_g1580B (.Q(g1580B),.SE(test_seB),.SI(g369B),.D(g6500B),.CK(CKB));
SDFF_X1 U_g1736B (.Q(g1736B),.SE(test_seB),.SI(g1580B),.D(g5392B),.CK(CKB));
SDFF_X1 U_g39B (.Q(g39B),.SE(test_seB),.SI(g1736B),.D(g10663B),.CK(CKB));
SDFF_X1 U_g1651B (.Q(g1651B),.SE(test_seB),.SI(g39B),.D(g10782B),.CK(CKB));
SDFF_X1 U_g1424B (.Q(g1424B),.SE(test_seB),.SI(g1651B),.D(g6216B),.CK(CKB));
SDFF_X1 U_g1737B (.Q(g1737B),.SE(test_seB),.SI(g1424B),.D(g1736B),.CK(CKB));
SDFF_X1 U_g1672B (.Q(g1672B),.SE(test_seB),.SI(g1737B),.D(g10858B),.CK(CKB));
SDFF_X1 U_g1077B (.Q(g1077B),.SE(test_seB),.SI(g1672B),.D(g5914B),.CK(CKB));
SDFF_X1 U_g1231B (.Q(g1231B),.SE(test_seB),.SI(g1077B),.D(g7590B),.CK(CKB));
SDFF_X1 U_g4B (.Q(g4B),.SE(test_seB),.SI(g1231B),.D(g6656B),.CK(CKB));
SDFF_X1 U_g774B (.Q(g774B),.SE(test_seB),.SI(g4B),.D(g6728B),.CK(CKB));
SDFF_X1 U_g1104B (.Q(g1104B),.SE(test_seB),.SI(g774B),.D(g5126B),.CK(CKB));
SDFF_X1 U_g1304B (.Q(g1304B),.SE(test_seB),.SI(g1104B),.D(g7290B),.CK(CKB));
SDFF_X1 U_g243B (.Q(g243B),.SE(test_seB),.SI(g1304B),.D(g6841B),.CK(CKB));
SDFF_X1 U_g1499B (.Q(g1499B),.SE(test_seB),.SI(g243B),.D(g8041B),.CK(CKB));
SDFF_X1 U_g1044B (.Q(g1044B),.SE(test_seB),.SI(g1499B),.D(g7106B),.CK(CKB));
SDFF_X1 U_g1444B (.Q(g1444B),.SE(test_seB),.SI(g1044B),.D(g8766B),.CK(CKB));
SDFF_X1 U_g757B (.Q(g757B),.SE(test_seB),.SI(g1444B),.D(g10788B),.CK(CKB));
SDFF_X1 U_g786B (.Q(g786B),.SE(test_seB),.SI(g757B),.D(g8019B),.CK(CKB));
SDFF_X1 U_g1543B (.Q(g1543B),.SE(test_seB),.SI(g786B),.D(g6545B),.CK(CKB));
SDFF_X1 U_g552B (.Q(g552B),.SE(test_seB),.SI(g1543B),.D(g10856B),.CK(CKB));
SDFF_X1 U_g315B (.Q(g315B),.SE(test_seB),.SI(g552B),.D(g256B),.CK(CKB));
SDFF_X1 U_g1534B (.Q(g1534B),.SE(test_seB),.SI(g315B),.D(g6533B),.CK(CKB));
SDFF_X1 U_g622B (.Q(g622B),.SE(test_seB),.SI(g1534B),.D(g8820B),.CK(CKB));
SDFF_X1 U_g1927B (.Q(g1927B),.SE(test_seB),.SI(g622B),.D(g8941B),.CK(CKB));
SDFF_X1 U_g1660B (.Q(g1660B),.SE(test_seB),.SI(g1927B),.D(g10859B),.CK(CKB));
SDFF_X1 U_g278B (.Q(g278B),.SE(test_seB),.SI(g1660B),.D(g6922B),.CK(CKB));
SDFF_X1 U_g1436B (.Q(g1436B),.SE(test_seB),.SI(g278B),.D(g8772B),.CK(CKB));
SDFF_X1 U_g718B (.Q(g718B),.SE(test_seB),.SI(g1436B),.D(g8433B),.CK(CKB));
SDFF_X1 U_g76B (.Q(g76B),.SE(test_seB),.SI(g718B),.D(g6526B),.CK(CKB));
SDFF_X1 U_g554B (.Q(g554B),.SE(test_seB),.SI(g76B),.D(g10793B),.CK(CKB));
SDFF_X1 U_g496B (.Q(g496B),.SE(test_seB),.SI(g554B),.D(g11333B),.CK(CKB));
SDFF_X1 U_g981B (.Q(g981B),.SE(test_seB),.SI(g496B),.D(g11392B),.CK(CKB));
SDFF_X1 U_g878B (.Q(g878B),.SE(test_seB),.SI(g981B),.D(g3506B),.CK(CKB));
SDFF_X1 U_g590B (.Q(g590B),.SE(test_seB),.SI(g878B),.D(g1713B),.CK(CKB));
SDFF_X1 U_g829B (.Q(g829B),.SE(test_seB),.SI(g590B),.D(g794B),.CK(CKB));
SDFF_X1 U_g1095B (.Q(g1095B),.SE(test_seB),.SI(g829B),.D(g6093B),.CK(CKB));
SDFF_X1 U_g704B (.Q(g704B),.SE(test_seB),.SI(g1095B),.D(g8889B),.CK(CKB));
SDFF_X1 U_g1265B (.Q(g1265B),.SE(test_seB),.SI(g704B),.D(g7302B),.CK(CKB));
SDFF_X1 U_g1786B (.Q(g1786B),.SE(test_seB),.SI(g1265B),.D(g6525B),.CK(CKB));
SDFF_X1 U_g682B (.Q(g682B),.SE(test_seB),.SI(g1786B),.D(g8429B),.CK(CKB));
SDFF_X1 U_g1296B (.Q(g1296B),.SE(test_seB),.SI(g682B),.D(g7292B),.CK(CKB));
SDFF_X1 U_g587B (.Q(g587B),.SE(test_seB),.SI(g1296B),.D(g104B),.CK(CKB));
SDFF_X1 U_g52B (.Q(g52B),.SE(test_seB),.SI(g587B),.D(g6621B),.CK(CKB));
SDFF_X1 U_g646B (.Q(g646B),.SE(test_seB),.SI(g52B),.D(g7134B),.CK(CKB));
SDFF_X1 U_g327B (.Q(g327B),.SE(test_seB),.SI(g646B),.D(g260B),.CK(CKB));
SDFF_X1 U_g1389B (.Q(g1389B),.SE(test_seB),.SI(g327B),.D(g6333B),.CK(CKB));
SDFF_X1 U_g1371B (.Q(g1371B),.SE(test_seB),.SI(g1389B),.D(g6826B),.CK(CKB));
SDFF_X1 U_g1956B (.Q(g1956B),.SE(test_seB),.SI(g1371B),.D(g1955B),.CK(CKB));
SDFF_X1 U_g1675B (.Q(g1675B),.SE(test_seB),.SI(g1956B),.D(g10860B),.CK(CKB));
SDFF_X1 U_g354B (.Q(g354B),.SE(test_seB),.SI(g1675B),.D(g11483B),.CK(CKB));
SDFF_X1 U_g113B (.Q(g113B),.SE(test_seB),.SI(g354B),.D(g6392B),.CK(CKB));
SDFF_X1 U_g639B (.Q(g639B),.SE(test_seB),.SI(g113B),.D(g7626B),.CK(CKB));
SDFF_X1 U_g1684B (.Q(g1684B),.SE(test_seB),.SI(g639B),.D(g10866B),.CK(CKB));
SDFF_X1 U_g1639B (.Q(g1639B),.SE(test_seB),.SI(g1684B),.D(g8193B),.CK(CKB));
SDFF_X1 U_g1791B (.Q(g1791B),.SE(test_seB),.SI(g1639B),.D(g6983B),.CK(CKB));
SDFF_X1 U_g248B (.Q(g248B),.SE(test_seB),.SI(g1791B),.D(g6839B),.CK(CKB));
SDFF_X1 U_g1707B (.Q(g1707B),.SE(test_seB),.SI(g248B),.D(g4076B),.CK(CKB));
SDFF_X1 U_g1759B (.Q(g1759B),.SE(test_seB),.SI(g1707B),.D(g4293B),.CK(CKB));
SDFF_X1 U_g351B (.Q(g351B),.SE(test_seB),.SI(g1759B),.D(g11482B),.CK(CKB));
SDFF_X1 U_g1957B (.Q(g1957B),.SE(test_seB),.SI(g351B),.D(g1956B),.CK(CKB));
SDFF_X1 U_g1604B (.Q(g1604B),.SE(test_seB),.SI(g1957B),.D(g6507B),.CK(CKB));
SDFF_X1 U_g1098B (.Q(g1098B),.SE(test_seB),.SI(g1604B),.D(g6096B),.CK(CKB));
SDFF_X1 U_g932B (.Q(g932B),.SE(test_seB),.SI(g1098B),.D(g8250B),.CK(CKB));
SDFF_X1 U_g126B (.Q(g126B),.SE(test_seB),.SI(g932B),.D(I8503B),.CK(CKB));
SDFF_X1 U_g1896B (.Q(g1896B),.SE(test_seB),.SI(g126B),.D(g8282B),.CK(CKB));
SDFF_X1 U_g736B (.Q(g736B),.SE(test_seB),.SI(g1896B),.D(g8435B),.CK(CKB));
SDFF_X1 U_g1019B (.Q(g1019B),.SE(test_seB),.SI(g736B),.D(g6924B),.CK(CKB));
SDFF_X1 U_g1362B (.Q(g1362B),.SE(test_seB),.SI(g1019B),.D(g6819B),.CK(CKB));
SDFF_X1 U_g745B (.Q(g745B),.SE(test_seB),.SI(g1362B),.D(g746B),.CK(CKB));
SDFF_X1 U_g1419B (.Q(g1419B),.SE(test_seB),.SI(g745B),.D(g6244B),.CK(CKB));
SDFF_X1 U_g58B (.Q(g58B),.SE(test_seB),.SI(g1419B),.D(g6627B),.CK(CKB));
SDFF_X1 U_g32B (.Q(g32B),.SE(test_seB),.SI(g58B),.D(g11286B),.CK(CKB));
SDFF_X1 U_g876B (.Q(g876B),.SE(test_seB),.SI(g32B),.D(g878B),.CK(CKB));
SDFF_X1 U_g1086B (.Q(g1086B),.SE(test_seB),.SI(g876B),.D(g6071B),.CK(CKB));
SDFF_X1 U_g1486B (.Q(g1486B),.SE(test_seB),.SI(g1086B),.D(g8046B),.CK(CKB));
SDFF_X1 U_g1730B (.Q(g1730B),.SE(test_seB),.SI(g1486B),.D(g10707B),.CK(CKB));
SDFF_X1 U_g1504B (.Q(g1504B),.SE(test_seB),.SI(g1730B),.D(g6198B),.CK(CKB));
SDFF_X1 U_g1470B (.Q(g1470B),.SE(test_seB),.SI(g1504B),.D(g8051B),.CK(CKB));
SDFF_X1 U_g822B (.Q(g822B),.SE(test_seB),.SI(g1470B),.D(g8024B),.CK(CKB));
SDFF_X1 U_g583B (.Q(g583B),.SE(test_seB),.SI(g822B),.D(g29B),.CK(CKB));
SDFF_X1 U_g1678B (.Q(g1678B),.SE(test_seB),.SI(g583B),.D(g10862B),.CK(CKB));
SDFF_X1 U_g174B (.Q(g174B),.SE(test_seB),.SI(g1678B),.D(g8050B),.CK(CKB));
SDFF_X1 U_g1766B (.Q(g1766B),.SE(test_seB),.SI(g174B),.D(g7133B),.CK(CKB));
SDFF_X1 U_g1801B (.Q(g1801B),.SE(test_seB),.SI(g1766B),.D(g7930B),.CK(CKB));
SDFF_X1 U_g186B (.Q(g186B),.SE(test_seB),.SI(g1801B),.D(g6832B),.CK(CKB));
SDFF_X1 U_g959B (.Q(g959B),.SE(test_seB),.SI(g186B),.D(g11308B),.CK(CKB));
SDFF_X1 U_g1169B (.Q(g1169B),.SE(test_seB),.SI(g959B),.D(g5189B),.CK(CKB));
SDFF_X1 U_g1007B (.Q(g1007B),.SE(test_seB),.SI(g1169B),.D(g6918B),.CK(CKB));
SDFF_X1 U_g1407B (.Q(g1407B),.SE(test_seB),.SI(g1007B),.D(g8769B),.CK(CKB));
SDFF_X1 U_g1059B (.Q(g1059B),.SE(test_seB),.SI(g1407B),.D(g7236B),.CK(CKB));
SDFF_X1 U_g1868B (.Q(g1868B),.SE(test_seB),.SI(g1059B),.D(g6909B),.CK(CKB));
SDFF_X1 U_g758B (.Q(g758B),.SE(test_seB),.SI(g1868B),.D(g4940B),.CK(CKB));
SDFF_X1 U_g1718B (.Q(g1718B),.SE(test_seB),.SI(g758B),.D(g5404B),.CK(CKB));
SDFF_X1 U_g396B (.Q(g396B),.SE(test_seB),.SI(g1718B),.D(g11265B),.CK(CKB));
SDFF_X1 U_g1015B (.Q(g1015B),.SE(test_seB),.SI(g396B),.D(g6930B),.CK(CKB));
SDFF_X1 U_g38B (.Q(g38B),.SE(test_seB),.SI(g1015B),.D(g10726B),.CK(CKB));
SDFF_X1 U_g632B (.Q(g632B),.SE(test_seB),.SI(g38B),.D(g4891B),.CK(CKB));
SDFF_X1 U_g1415B (.Q(g1415B),.SE(test_seB),.SI(g632B),.D(g6224B),.CK(CKB));
SDFF_X1 U_g1227B (.Q(g1227B),.SE(test_seB),.SI(g1415B),.D(g7586B),.CK(CKB));
SDFF_X1 U_g1721B (.Q(g1721B),.SE(test_seB),.SI(g1227B),.D(g10770B),.CK(CKB));
SDFF_X1 U_g882B (.Q(g882B),.SE(test_seB),.SI(g1721B),.D(g883B),.CK(CKB));
SDFF_X1 U_g16B (.Q(g16B),.SE(test_seB),.SI(g882B),.D(g3524B),.CK(CKB));
SDFF_X1 U_g284B (.Q(g284B),.SE(test_seB),.SI(g16B),.D(g6934B),.CK(CKB));
SDFF_X1 U_g426B (.Q(g426B),.SE(test_seB),.SI(g284B),.D(g11256B),.CK(CKB));
SDFF_X1 U_g219B (.Q(g219B),.SE(test_seB),.SI(g426B),.D(g6824B),.CK(CKB));
SDFF_X1 U_g1216B (.Q(g1216B),.SE(test_seB),.SI(g219B),.D(g1360B),.CK(CKB));
SDFF_X1 U_g806B (.Q(g806B),.SE(test_seB),.SI(g1216B),.D(g6126B),.CK(CKB));
SDFF_X1 U_g1428B (.Q(g1428B),.SE(test_seB),.SI(g806B),.D(g8767B),.CK(CKB));
SDFF_X1 U_g579B (.Q(g579B),.SE(test_seB),.SI(g1428B),.D(g102B),.CK(CKB));
SDFF_X1 U_g1564B (.Q(g1564B),.SE(test_seB),.SI(g579B),.D(g6546B),.CK(CKB));
SDFF_X1 U_g1741B (.Q(g1741B),.SE(test_seB),.SI(g1564B),.D(g4238B),.CK(CKB));
SDFF_X1 U_g225B (.Q(g225B),.SE(test_seB),.SI(g1741B),.D(g6823B),.CK(CKB));
SDFF_X1 U_g281B (.Q(g281B),.SE(test_seB),.SI(g225B),.D(g6928B),.CK(CKB));
SDFF_X1 U_g1308B (.Q(g1308B),.SE(test_seB),.SI(g281B),.D(g11602B),.CK(CKB));
SDFF_X1 U_g611B (.Q(g611B),.SE(test_seB),.SI(g1308B),.D(g9721B),.CK(CKB));
SDFF_X1 U_g631B (.Q(g631B),.SE(test_seB),.SI(g611B),.D(g4890B),.CK(CKB));
SDFF_X1 U_g1217B (.Q(g1217B),.SE(test_seB),.SI(g631B),.D(g9525B),.CK(CKB));
SDFF_X1 U_g1589B (.Q(g1589B),.SE(test_seB),.SI(g1217B),.D(g6524B),.CK(CKB));
SDFF_X1 U_g1466B (.Q(g1466B),.SE(test_seB),.SI(g1589B),.D(g8045B),.CK(CKB));
SDFF_X1 U_g1571B (.Q(g1571B),.SE(test_seB),.SI(g1466B),.D(g6469B),.CK(CKB));
SDFF_X1 U_g1861B (.Q(g1861B),.SE(test_seB),.SI(g1571B),.D(g6471B),.CK(CKB));
SDFF_X1 U_g1365B (.Q(g1365B),.SE(test_seB),.SI(g1861B),.D(g6821B),.CK(CKB));
SDFF_X1 U_g1448B (.Q(g1448B),.SE(test_seB),.SI(g1365B),.D(g11514B),.CK(CKB));
SDFF_X1 U_g1711B (.Q(g1711B),.SE(test_seB),.SI(g1448B),.D(g5403B),.CK(CKB));
SDFF_X1 U_g1133B (.Q(g1133B),.SE(test_seB),.SI(g1711B),.D(g4480B),.CK(CKB));
SDFF_X1 U_g1333B (.Q(g1333B),.SE(test_seB),.SI(g1133B),.D(g11610B),.CK(CKB));
SDFF_X1 U_g153B (.Q(g153B),.SE(test_seB),.SI(g1333B),.D(g7843B),.CK(CKB));
SDFF_X1 U_g962B (.Q(g962B),.SE(test_seB),.SI(g153B),.D(g11310B),.CK(CKB));
SDFF_X1 U_g766B (.Q(g766B),.SE(test_seB),.SI(g962B),.D(g5536B),.CK(CKB));
SDFF_X1 U_g588B (.Q(g588B),.SE(test_seB),.SI(g766B),.D(g28B),.CK(CKB));
SDFF_X1 U_g486B (.Q(g486B),.SE(test_seB),.SI(g588B),.D(g11331B),.CK(CKB));
SDFF_X1 U_g471B (.Q(g471B),.SE(test_seB),.SI(g486B),.D(g11380B),.CK(CKB));
SDFF_X1 U_g1397B (.Q(g1397B),.SE(test_seB),.SI(g471B),.D(g6838B),.CK(CKB));
SDFF_X1 U_g580B (.Q(g580B),.SE(test_seB),.SI(g1397B),.D(g103B),.CK(CKB));
SDFF_X1 U_g1950B (.Q(g1950B),.SE(test_seB),.SI(g580B),.D(g8288B),.CK(CKB));
SDFF_X1 U_g756B (.Q(g756B),.SE(test_seB),.SI(g1950B),.D(g755B),.CK(CKB));
SDFF_X1 U_g635B (.Q(g635B),.SE(test_seB),.SI(g756B),.D(g4892B),.CK(CKB));
SDFF_X1 U_g1101B (.Q(g1101B),.SE(test_seB),.SI(g635B),.D(g5390B),.CK(CKB));
SDFF_X1 U_g549B (.Q(g549B),.SE(test_seB),.SI(g1101B),.D(g10855B),.CK(CKB));
SDFF_X1 U_g1041B (.Q(g1041B),.SE(test_seB),.SI(g549B),.D(g7258B),.CK(CKB));
SDFF_X1 U_g105B (.Q(g105B),.SE(test_seB),.SI(g1041B),.D(g10898B),.CK(CKB));
SDFF_X1 U_g1669B (.Q(g1669B),.SE(test_seB),.SI(g105B),.D(g10865B),.CK(CKB));
SDFF_X1 U_g1368B (.Q(g1368B),.SE(test_seB),.SI(g1669B),.D(g6822B),.CK(CKB));
SDFF_X1 U_g1531B (.Q(g1531B),.SE(test_seB),.SI(g1368B),.D(g6528B),.CK(CKB));
SDFF_X1 U_g1458B (.Q(g1458B),.SE(test_seB),.SI(g1531B),.D(g6180B),.CK(CKB));
SDFF_X1 U_g572B (.Q(g572B),.SE(test_seB),.SI(g1458B),.D(g10718B),.CK(CKB));
SDFF_X1 U_g1011B (.Q(g1011B),.SE(test_seB),.SI(g572B),.D(g6912B),.CK(CKB));
SDFF_X1 U_g33B (.Q(g33B),.SE(test_seB),.SI(g1011B),.D(g10719B),.CK(CKB));
SDFF_X1 U_g1411B (.Q(g1411B),.SE(test_seB),.SI(g33B),.D(g6234B),.CK(CKB));
SDFF_X1 U_g1074B (.Q(g1074B),.SE(test_seB),.SI(g1411B),.D(g6099B),.CK(CKB));
SDFF_X1 U_g444B (.Q(g444B),.SE(test_seB),.SI(g1074B),.D(g11259B),.CK(CKB));
SDFF_X1 U_g1474B (.Q(g1474B),.SE(test_seB),.SI(g444B),.D(g8039B),.CK(CKB));
SDFF_X1 U_g1080B (.Q(g1080B),.SE(test_seB),.SI(g1474B),.D(g6059B),.CK(CKB));
SDFF_X1 U_g1713B (.Q(g1713B),.SE(test_seB),.SI(g1080B),.D(g5396B),.CK(CKB));
SDFF_X1 U_g333B (.Q(g333B),.SE(test_seB),.SI(g1713B),.D(g262B),.CK(CKB));
SDFF_X1 U_g269B (.Q(g269B),.SE(test_seB),.SI(g333B),.D(g6906B),.CK(CKB));
SDFF_X1 U_g401B (.Q(g401B),.SE(test_seB),.SI(g269B),.D(g11266B),.CK(CKB));
SDFF_X1 U_g1857B (.Q(g1857B),.SE(test_seB),.SI(g401B),.D(g11294B),.CK(CKB));
SDFF_X1 U_g9B (.Q(g9B),.SE(test_seB),.SI(g1857B),.D(g5421B),.CK(CKB));
SDFF_X1 U_g664B (.Q(g664B),.SE(test_seB),.SI(g9B),.D(g8649B),.CK(CKB));
SDFF_X1 U_g965B (.Q(g965B),.SE(test_seB),.SI(g664B),.D(g11312B),.CK(CKB));
SDFF_X1 U_g1400B (.Q(g1400B),.SE(test_seB),.SI(g965B),.D(g6840B),.CK(CKB));
SDFF_X1 U_g309B (.Q(g309B),.SE(test_seB),.SI(g1400B),.D(g254B),.CK(CKB));
SDFF_X1 U_g814B (.Q(g814B),.SE(test_seB),.SI(g309B),.D(g7202B),.CK(CKB));
SDFF_X1 U_g231B (.Q(g231B),.SE(test_seB),.SI(g814B),.D(g6834B),.CK(CKB));
SDFF_X1 U_g557B (.Q(g557B),.SE(test_seB),.SI(g231B),.D(g10795B),.CK(CKB));
SDFF_X1 U_g586B (.Q(g586B),.SE(test_seB),.SI(g557B),.D(g103B),.CK(CKB));
SDFF_X1 U_g869B (.Q(g869B),.SE(test_seB),.SI(g586B),.D(g875B),.CK(CKB));
SDFF_X1 U_g1383B (.Q(g1383B),.SE(test_seB),.SI(g869B),.D(g6831B),.CK(CKB));
SDFF_X1 U_g158B (.Q(g158B),.SE(test_seB),.SI(g1383B),.D(g8060B),.CK(CKB));
SDFF_X1 U_g627B (.Q(g627B),.SE(test_seB),.SI(g158B),.D(g4893B),.CK(CKB));
SDFF_X1 U_g1023B (.Q(g1023B),.SE(test_seB),.SI(g627B),.D(g7244B),.CK(CKB));
SDFF_X1 U_g259B (.Q(g259B),.SE(test_seB),.SI(g1023B),.D(g6026B),.CK(CKB));
SDFF_X1 U_g1361B (.Q(g1361B),.SE(test_seB),.SI(g259B),.D(g1206B),.CK(CKB));
SDFF_X1 U_g1327B (.Q(g1327B),.SE(test_seB),.SI(g1361B),.D(g11608B),.CK(CKB));
SDFF_X1 U_g654B (.Q(g654B),.SE(test_seB),.SI(g1327B),.D(g7660B),.CK(CKB));
SDFF_X1 U_g293B (.Q(g293B),.SE(test_seB),.SI(g654B),.D(g6911B),.CK(CKB));
SDFF_X1 U_g1346B (.Q(g1346B),.SE(test_seB),.SI(g293B),.D(g11640B),.CK(CKB));
SDFF_X1 U_g1633B (.Q(g1633B),.SE(test_seB),.SI(g1346B),.D(g8777B),.CK(CKB));
SDFF_X1 U_g1753B (.Q(g1753B),.SE(test_seB),.SI(g1633B),.D(g4274B),.CK(CKB));
SDFF_X1 U_g1508B (.Q(g1508B),.SE(test_seB),.SI(g1753B),.D(g6215B),.CK(CKB));
SDFF_X1 U_g1240B (.Q(g1240B),.SE(test_seB),.SI(g1508B),.D(g7297B),.CK(CKB));
SDFF_X1 U_g538B (.Q(g538B),.SE(test_seB),.SI(g1240B),.D(g11326B),.CK(CKB));
SDFF_X1 U_g416B (.Q(g416B),.SE(test_seB),.SI(g538B),.D(g11269B),.CK(CKB));
SDFF_X1 U_g542B (.Q(g542B),.SE(test_seB),.SI(g416B),.D(g11325B),.CK(CKB));
SDFF_X1 U_g1681B (.Q(g1681B),.SE(test_seB),.SI(g542B),.D(g10864B),.CK(CKB));
SDFF_X1 U_g374B (.Q(g374B),.SE(test_seB),.SI(g1681B),.D(g11290B),.CK(CKB));
SDFF_X1 U_g563B (.Q(g563B),.SE(test_seB),.SI(g374B),.D(g10798B),.CK(CKB));
SDFF_X1 U_g1914B (.Q(g1914B),.SE(test_seB),.SI(g563B),.D(g8284B),.CK(CKB));
SDFF_X1 U_g530B (.Q(g530B),.SE(test_seB),.SI(g1914B),.D(g11328B),.CK(CKB));
SDFF_X1 U_g575B (.Q(g575B),.SE(test_seB),.SI(g530B),.D(g10800B),.CK(CKB));
SDFF_X1 U_g1936B (.Q(g1936B),.SE(test_seB),.SI(g575B),.D(g8944B),.CK(CKB));
SDFF_X1 U_g55B (.Q(g55B),.SE(test_seB),.SI(g1936B),.D(g7183B),.CK(CKB));
SDFF_X1 U_g1117B (.Q(g1117B),.SE(test_seB),.SI(g55B),.D(g4465B),.CK(CKB));
SDFF_X1 U_g1317B (.Q(g1317B),.SE(test_seB),.SI(g1117B),.D(g1356B),.CK(CKB));
SDFF_X1 U_g357B (.Q(g357B),.SE(test_seB),.SI(g1317B),.D(g11484B),.CK(CKB));
SDFF_X1 U_g386B (.Q(g386B),.SE(test_seB),.SI(g357B),.D(g11263B),.CK(CKB));
SDFF_X1 U_g1601B (.Q(g1601B),.SE(test_seB),.SI(g386B),.D(g6501B),.CK(CKB));
SDFF_X1 U_g553B (.Q(g553B),.SE(test_seB),.SI(g1601B),.D(g10857B),.CK(CKB));
SDFF_X1 U_g166B (.Q(g166B),.SE(test_seB),.SI(g553B),.D(g6757B),.CK(CKB));
SDFF_X1 U_g501B (.Q(g501B),.SE(test_seB),.SI(g166B),.D(g11334B),.CK(CKB));
SDFF_X1 U_g262B (.Q(g262B),.SE(test_seB),.SI(g501B),.D(g6042B),.CK(CKB));
SDFF_X1 U_g1840B (.Q(g1840B),.SE(test_seB),.SI(g262B),.D(g8384B),.CK(CKB));
SDFF_X1 U_g70B (.Q(g70B),.SE(test_seB),.SI(g1840B),.D(g6653B),.CK(CKB));
SDFF_X1 U_g318B (.Q(g318B),.SE(test_seB),.SI(g70B),.D(g257B),.CK(CKB));
SDFF_X1 U_g1356B (.Q(g1356B),.SE(test_seB),.SI(g318B),.D(g5763B),.CK(CKB));
SDFF_X1 U_g794B (.Q(g794B),.SE(test_seB),.SI(g1356B),.D(g5849B),.CK(CKB));
SDFF_X1 U_g36B (.Q(g36B),.SE(test_seB),.SI(g794B),.D(g10722B),.CK(CKB));
SDFF_X1 U_g302B (.Q(g302B),.SE(test_seB),.SI(g36B),.D(g6929B),.CK(CKB));
SDFF_X1 U_g342B (.Q(g342B),.SE(test_seB),.SI(g302B),.D(g11488B),.CK(CKB));
SDFF_X1 U_g1250B (.Q(g1250B),.SE(test_seB),.SI(g342B),.D(g7299B),.CK(CKB));
SDFF_X1 U_g1163B (.Q(g1163B),.SE(test_seB),.SI(g1250B),.D(g4330B),.CK(CKB));
SDFF_X1 U_g1810B (.Q(g1810B),.SE(test_seB),.SI(g1163B),.D(g1958B),.CK(CKB));
SDFF_X1 U_g1032B (.Q(g1032B),.SE(test_seB),.SI(g1810B),.D(g7257B),.CK(CKB));
SDFF_X1 U_g1432B (.Q(g1432B),.SE(test_seB),.SI(g1032B),.D(g8775B),.CK(CKB));
SDFF_X1 U_g1053B (.Q(g1053B),.SE(test_seB),.SI(g1432B),.D(g7225B),.CK(CKB));
SDFF_X1 U_g1453B (.Q(g1453B),.SE(test_seB),.SI(g1053B),.D(g5770B),.CK(CKB));
SDFF_X1 U_g363B (.Q(g363B),.SE(test_seB),.SI(g1453B),.D(g11486B),.CK(CKB));
SDFF_X1 U_g330B (.Q(g330B),.SE(test_seB),.SI(g363B),.D(g261B),.CK(CKB));
SDFF_X1 U_g1157B (.Q(g1157B),.SE(test_seB),.SI(g330B),.D(g4338B),.CK(CKB));
SDFF_X1 U_g1357B (.Q(g1357B),.SE(test_seB),.SI(g1157B),.D(g4500B),.CK(CKB));
SDFF_X1 U_g35B (.Q(g35B),.SE(test_seB),.SI(g1357B),.D(g10721B),.CK(CKB));
SDFF_X1 U_g928B (.Q(g928B),.SE(test_seB),.SI(g35B),.D(g8147B),.CK(CKB));
SDFF_X1 U_g261B (.Q(g261B),.SE(test_seB),.SI(g928B),.D(g6038B),.CK(CKB));
SDFF_X1 U_g516B (.Q(g516B),.SE(test_seB),.SI(g261B),.D(g11337B),.CK(CKB));
SDFF_X1 U_g254B (.Q(g254B),.SE(test_seB),.SI(g516B),.D(g6045B),.CK(CKB));
SDFF_X1 U_g778B (.Q(g778B),.SE(test_seB),.SI(g254B),.D(g7191B),.CK(CKB));
SDFF_X1 U_g861B (.Q(g861B),.SE(test_seB),.SI(g778B),.D(g826B),.CK(CKB));
SDFF_X1 U_g1627B (.Q(g1627B),.SE(test_seB),.SI(g861B),.D(g8774B),.CK(CKB));
SDFF_X1 U_g1292B (.Q(g1292B),.SE(test_seB),.SI(g1627B),.D(g7293B),.CK(CKB));
SDFF_X1 U_g290B (.Q(g290B),.SE(test_seB),.SI(g1292B),.D(g6907B),.CK(CKB));
SDFF_X1 U_g1850B (.Q(g1850B),.SE(test_seB),.SI(g290B),.D(g4903B),.CK(CKB));
SDFF_X1 U_g770B (.Q(g770B),.SE(test_seB),.SI(g1850B),.D(g6123B),.CK(CKB));
SDFF_X1 U_g1583B (.Q(g1583B),.SE(test_seB),.SI(g770B),.D(g6506B),.CK(CKB));
SDFF_X1 U_g466B (.Q(g466B),.SE(test_seB),.SI(g1583B),.D(g11376B),.CK(CKB));
SDFF_X1 U_g1561B (.Q(g1561B),.SE(test_seB),.SI(g466B),.D(g6542B),.CK(CKB));
SDFF_X1 U_g1527B (.Q(g1527B),.SE(test_seB),.SI(g1561B),.D(I8503B),.CK(CKB));
SDFF_X1 U_g1546B (.Q(g1546B),.SE(test_seB),.SI(g1527B),.D(g6551B),.CK(CKB));
SDFF_X1 U_g287B (.Q(g287B),.SE(test_seB),.SI(g1546B),.D(g6901B),.CK(CKB));
SDFF_X1 U_g560B (.Q(g560B),.SE(test_seB),.SI(g287B),.D(g10797B),.CK(CKB));
SDFF_X1 U_g617B (.Q(g617B),.SE(test_seB),.SI(g560B),.D(g8505B),.CK(CKB));
SDFF_X1 U_g17B (.Q(g17B),.SE(test_seB),.SI(g617B),.D(g4117B),.CK(CKB));
SDFF_X1 U_g336B (.Q(g336B),.SE(test_seB),.SI(g17B),.D(g11647B),.CK(CKB));
SDFF_X1 U_g456B (.Q(g456B),.SE(test_seB),.SI(g336B),.D(g11340B),.CK(CKB));
SDFF_X1 U_g305B (.Q(g305B),.SE(test_seB),.SI(g456B),.D(g253B),.CK(CKB));
SDFF_X1 U_g345B (.Q(g345B),.SE(test_seB),.SI(g305B),.D(g11625B),.CK(CKB));
SDFF_X1 U_g8B (.Q(g8B),.SE(test_seB),.SI(g345B),.D(g636B),.CK(CKB));
SDFF_X1 U_g1771B (.Q(g1771B),.SE(test_seB),.SI(g8B),.D(g6502B),.CK(CKB));
SDFF_X1 U_g865B (.Q(g865B),.SE(test_seB),.SI(g1771B),.D(g7981B),.CK(CKB));
SDFF_X1 U_g255B (.Q(g255B),.SE(test_seB),.SI(g865B),.D(g6049B),.CK(CKB));
SDFF_X1 U_g1945B (.Q(g1945B),.SE(test_seB),.SI(g255B),.D(g8945B),.CK(CKB));
SDFF_X1 U_g1738B (.Q(g1738B),.SE(test_seB),.SI(g1945B),.D(g4231B),.CK(CKB));
SDFF_X1 U_g1478B (.Q(g1478B),.SE(test_seB),.SI(g1738B),.D(g8040B),.CK(CKB));
SDFF_X1 U_g1035B (.Q(g1035B),.SE(test_seB),.SI(g1478B),.D(g7203B),.CK(CKB));
SDFF_X1 U_g1959B (.Q(g1959B),.SE(test_seB),.SI(g1035B),.D(I5254B),.CK(CKB));
SDFF_X1 U_g1690B (.Q(g1690B),.SE(test_seB),.SI(g1959B),.D(g6155B),.CK(CKB));
SDFF_X1 U_g1482B (.Q(g1482B),.SE(test_seB),.SI(g1690B),.D(g8043B),.CK(CKB));
SDFF_X1 U_g1110B (.Q(g1110B),.SE(test_seB),.SI(g1482B),.D(g5173B),.CK(CKB));
SDFF_X1 U_g296B (.Q(g296B),.SE(test_seB),.SI(g1110B),.D(g6916B),.CK(CKB));
SDFF_X1 U_g1663B (.Q(g1663B),.SE(test_seB),.SI(g296B),.D(g10861B),.CK(CKB));
SDFF_X1 U_g700B (.Q(g700B),.SE(test_seB),.SI(g1663B),.D(g8431B),.CK(CKB));
SDFF_X1 U_g1762B (.Q(g1762B),.SE(test_seB),.SI(g700B),.D(g4309B),.CK(CKB));
SDFF_X1 U_g360B (.Q(g360B),.SE(test_seB),.SI(g1762B),.D(g11485B),.CK(CKB));
SDFF_X1 U_g192B (.Q(g192B),.SE(test_seB),.SI(g360B),.D(g6334B),.CK(CKB));
SDFF_X1 U_g1657B (.Q(g1657B),.SE(test_seB),.SI(g192B),.D(g10767B),.CK(CKB));
SDFF_X1 U_g722B (.Q(g722B),.SE(test_seB),.SI(g1657B),.D(g8923B),.CK(CKB));
SDFF_X1 U_g61B (.Q(g61B),.SE(test_seB),.SI(g722B),.D(g7189B),.CK(CKB));
SDFF_X1 U_g566B (.Q(g566B),.SE(test_seB),.SI(g61B),.D(g10799B),.CK(CKB));
SDFF_X1 U_g1394B (.Q(g1394B),.SE(test_seB),.SI(g566B),.D(g6747B),.CK(CKB));
SDFF_X1 U_g1089B (.Q(g1089B),.SE(test_seB),.SI(g1394B),.D(g6080B),.CK(CKB));
SDFF_X1 U_g883B (.Q(g883B),.SE(test_seB),.SI(g1089B),.D(g3381B),.CK(CKB));
SDFF_X1 U_g1071B (.Q(g1071B),.SE(test_seB),.SI(g883B),.D(g5910B),.CK(CKB));
SDFF_X1 U_g986B (.Q(g986B),.SE(test_seB),.SI(g1071B),.D(g11393B),.CK(CKB));
SDFF_X1 U_g971B (.Q(g971B),.SE(test_seB),.SI(g986B),.D(g11349B),.CK(CKB));
SDFF_X1 U_g1955B (.Q(g1955B),.SE(test_seB),.SI(g971B),.D(g83B),.CK(CKB));
SDFF_X1 U_g143B (.Q(g143B),.SE(test_seB),.SI(g1955B),.D(g6439B),.CK(CKB));
SDFF_X1 U_g1814B (.Q(g1814B),.SE(test_seB),.SI(g143B),.D(g9266B),.CK(CKB));
SDFF_X1 U_g1038B (.Q(g1038B),.SE(test_seB),.SI(g1814B),.D(g7245B),.CK(CKB));
SDFF_X1 U_g1212B (.Q(g1212B),.SE(test_seB),.SI(g1038B),.D(g1217B),.CK(CKB));
SDFF_X1 U_g1918B (.Q(g1918B),.SE(test_seB),.SI(g1212B),.D(g8940B),.CK(CKB));
SDFF_X1 U_g782B (.Q(g782B),.SE(test_seB),.SI(g1918B),.D(g7705B),.CK(CKB));
SDFF_X1 U_g1822B (.Q(g1822B),.SE(test_seB),.SI(g782B),.D(g9269B),.CK(CKB));
SDFF_X1 U_g237B (.Q(g237B),.SE(test_seB),.SI(g1822B),.D(g6820B),.CK(CKB));
SDFF_X1 U_g746B (.Q(g746B),.SE(test_seB),.SI(g237B),.D(g756B),.CK(CKB));
SDFF_X1 U_g1062B (.Q(g1062B),.SE(test_seB),.SI(g746B),.D(g7240B),.CK(CKB));
SDFF_X1 U_g1462B (.Q(g1462B),.SE(test_seB),.SI(g1062B),.D(g8042B),.CK(CKB));
SDFF_X1 U_g178B (.Q(g178B),.SE(test_seB),.SI(g1462B),.D(g6759B),.CK(CKB));
SDFF_X1 U_g366B (.Q(g366B),.SE(test_seB),.SI(g178B),.D(g11487B),.CK(CKB));
SDFF_X1 U_g837B (.Q(g837B),.SE(test_seB),.SI(g366B),.D(g802B),.CK(CKB));
SDFF_X1 U_g599B (.Q(g599B),.SE(test_seB),.SI(g837B),.D(g9124B),.CK(CKB));
SDFF_X1 U_g1854B (.Q(g1854B),.SE(test_seB),.SI(g599B),.D(g11293B),.CK(CKB));
SDFF_X1 U_g944B (.Q(g944B),.SE(test_seB),.SI(g1854B),.D(g11298B),.CK(CKB));
SDFF_X1 U_g1941B (.Q(g1941B),.SE(test_seB),.SI(g944B),.D(g8287B),.CK(CKB));
SDFF_X1 U_g170B (.Q(g170B),.SE(test_seB),.SI(g1941B),.D(g8047B),.CK(CKB));
SDFF_X1 U_g1520B (.Q(g1520B),.SE(test_seB),.SI(g170B),.D(g6205B),.CK(CKB));
SDFF_X1 U_g686B (.Q(g686B),.SE(test_seB),.SI(g1520B),.D(g8885B),.CK(CKB));
SDFF_X1 U_g953B (.Q(g953B),.SE(test_seB),.SI(g686B),.D(g11305B),.CK(CKB));
SDFF_X1 U_g1958B (.Q(g1958B),.SE(test_seB),.SI(g953B),.D(g5556B),.CK(CKB));
SDFF_X1 U_g40B (.Q(g40B),.SE(test_seB),.SI(g1958B),.D(g10664B),.CK(CKB));
SDFF_X1 U_g1765B (.Q(g1765B),.SE(test_seB),.SI(g40B),.D(g2478B),.CK(CKB));
SDFF_X1 U_g1733B (.Q(g1733B),.SE(test_seB),.SI(g1765B),.D(g10711B),.CK(CKB));
SDFF_X1 U_g1270B (.Q(g1270B),.SE(test_seB),.SI(g1733B),.D(g7303B),.CK(CKB));
SDFF_X1 U_g1610B (.Q(g1610B),.SE(test_seB),.SI(g1270B),.D(g5194B),.CK(CKB));
SDFF_X1 U_g1796B (.Q(g1796B),.SE(test_seB),.SI(g1610B),.D(g7541B),.CK(CKB));
SDFF_X1 U_g1324B (.Q(g1324B),.SE(test_seB),.SI(g1796B),.D(g11607B),.CK(CKB));
SDFF_X1 U_g1540B (.Q(g1540B),.SE(test_seB),.SI(g1324B),.D(g6541B),.CK(CKB));
SDFF_X1 U_g1377B (.Q(g1377B),.SE(test_seB),.SI(g1540B),.D(g6827B),.CK(CKB));
SDFF_X1 U_g1206B (.Q(g1206B),.SE(test_seB),.SI(g1377B),.D(g4114B),.CK(CKB));
SDFF_X1 U_g491B (.Q(g491B),.SE(test_seB),.SI(g1206B),.D(g11332B),.CK(CKB));
SDFF_X1 U_g1849B (.Q(g1849B),.SE(test_seB),.SI(g491B),.D(g4902B),.CK(CKB));
SDFF_X1 U_g213B (.Q(g213B),.SE(test_seB),.SI(g1849B),.D(g6828B),.CK(CKB));
SDFF_X1 U_g1781B (.Q(g1781B),.SE(test_seB),.SI(g213B),.D(g6516B),.CK(CKB));
SDFF_X1 U_g1900B (.Q(g1900B),.SE(test_seB),.SI(g1781B),.D(g8938B),.CK(CKB));
SDFF_X1 U_g1245B (.Q(g1245B),.SE(test_seB),.SI(g1900B),.D(g7298B),.CK(CKB));
SDFF_X1 U_g108B (.Q(g108B),.SE(test_seB),.SI(g1245B),.D(g11561B),.CK(CKB));
SDFF_X1 U_g630B (.Q(g630B),.SE(test_seB),.SI(g108B),.D(g6672B),.CK(CKB));
SDFF_X1 U_g148B (.Q(g148B),.SE(test_seB),.SI(g630B),.D(g8048B),.CK(CKB));
SDFF_X1 U_g833B (.Q(g833B),.SE(test_seB),.SI(g148B),.D(g798B),.CK(CKB));
SDFF_X1 U_g1923B (.Q(g1923B),.SE(test_seB),.SI(g833B),.D(g8285B),.CK(CKB));
SDFF_X1 U_g936B (.Q(g936B),.SE(test_seB),.SI(g1923B),.D(g8254B),.CK(CKB));
SDFF_X1 U_g1215B (.Q(g1215B),.SE(test_seB),.SI(g936B),.D(g5229B),.CK(CKB));
SDFF_X1 U_g1314B (.Q(g1314B),.SE(test_seB),.SI(g1215B),.D(g11604B),.CK(CKB));
SDFF_X1 U_g849B (.Q(g849B),.SE(test_seB),.SI(g1314B),.D(g814B),.CK(CKB));
SDFF_X1 U_g1336B (.Q(g1336B),.SE(test_seB),.SI(g849B),.D(g11636B),.CK(CKB));
SDFF_X1 U_g272B (.Q(g272B),.SE(test_seB),.SI(g1336B),.D(g6910B),.CK(CKB));
SDFF_X1 U_g1806B (.Q(g1806B),.SE(test_seB),.SI(g272B),.D(g8173B),.CK(CKB));
SDFF_X1 U_g826B (.Q(g826B),.SE(test_seB),.SI(g1806B),.D(g8245B),.CK(CKB));
SDFF_X1 U_g1065B (.Q(g1065B),.SE(test_seB),.SI(g826B),.D(g7242B),.CK(CKB));
SDFF_X1 U_g1887B (.Q(g1887B),.SE(test_seB),.SI(g1065B),.D(g8281B),.CK(CKB));
SDFF_X1 U_g37B (.Q(g37B),.SE(test_seB),.SI(g1887B),.D(g10724B),.CK(CKB));
SDFF_X1 U_g968B (.Q(g968B),.SE(test_seB),.SI(g37B),.D(g11314B),.CK(CKB));
SDFF_X1 U_g1845B (.Q(g1845B),.SE(test_seB),.SI(g968B),.D(g4905B),.CK(CKB));
SDFF_X1 U_g1137B (.Q(g1137B),.SE(test_seB),.SI(g1845B),.D(g4484B),.CK(CKB));
SDFF_X1 U_g1891B (.Q(g1891B),.SE(test_seB),.SI(g1137B),.D(g8937B),.CK(CKB));
SDFF_X1 U_g1255B (.Q(g1255B),.SE(test_seB),.SI(g1891B),.D(g7300B),.CK(CKB));
SDFF_X1 U_g257B (.Q(g257B),.SE(test_seB),.SI(g1255B),.D(g6002B),.CK(CKB));
SDFF_X1 U_g874B (.Q(g874B),.SE(test_seB),.SI(g257B),.D(g9507B),.CK(CKB));
SDFF_X1 U_g591B (.Q(g591B),.SE(test_seB),.SI(g874B),.D(g9110B),.CK(CKB));
SDFF_X1 U_g731B (.Q(g731B),.SE(test_seB),.SI(g591B),.D(g8926B),.CK(CKB));
SDFF_X1 U_g636B (.Q(g636B),.SE(test_seB),.SI(g731B),.D(g8631B),.CK(CKB));
SDFF_X1 U_g1218B (.Q(g1218B),.SE(test_seB),.SI(g636B),.D(g7632B),.CK(CKB));
SDFF_X1 U_g605B (.Q(g605B),.SE(test_seB),.SI(g1218B),.D(g9150B),.CK(CKB));
SDFF_X1 U_g79B (.Q(g79B),.SE(test_seB),.SI(g605B),.D(g6531B),.CK(CKB));
SDFF_X1 U_g182B (.Q(g182B),.SE(test_seB),.SI(g79B),.D(g6786B),.CK(CKB));
SDFF_X1 U_g950B (.Q(g950B),.SE(test_seB),.SI(g182B),.D(g11303B),.CK(CKB));
SDFF_X1 U_g1129B (.Q(g1129B),.SE(test_seB),.SI(g950B),.D(g4477B),.CK(CKB));
SDFF_X1 U_g857B (.Q(g857B),.SE(test_seB),.SI(g1129B),.D(g822B),.CK(CKB));
SDFF_X1 U_g448B (.Q(g448B),.SE(test_seB),.SI(g857B),.D(g11258B),.CK(CKB));
SDFF_X1 U_g1828B (.Q(g1828B),.SE(test_seB),.SI(g448B),.D(g9272B),.CK(CKB));
SDFF_X1 U_g1727B (.Q(g1727B),.SE(test_seB),.SI(g1828B),.D(g10773B),.CK(CKB));
SDFF_X1 U_g1592B (.Q(g1592B),.SE(test_seB),.SI(g1727B),.D(g6470B),.CK(CKB));
SDFF_X1 U_g1703B (.Q(g1703B),.SE(test_seB),.SI(g1592B),.D(g5083B),.CK(CKB));
SDFF_X1 U_g1932B (.Q(g1932B),.SE(test_seB),.SI(g1703B),.D(g8286B),.CK(CKB));
SDFF_X1 U_g1624B (.Q(g1624B),.SE(test_seB),.SI(g1932B),.D(g8773B),.CK(CKB));
SDFF_X1 U_g26B (.Q(g26B),.SE(test_seB),.SI(g1624B),.D(g4158B),.CK(CKB));
SDFF_X1 U_g1068B (.Q(g1068B),.SE(test_seB),.SI(g26B),.D(g6054B),.CK(CKB));
SDFF_X1 U_g578B (.Q(g578B),.SE(test_seB),.SI(g1068B),.D(g101B),.CK(CKB));
SDFF_X1 U_g440B (.Q(g440B),.SE(test_seB),.SI(g578B),.D(g11260B),.CK(CKB));
SDFF_X1 U_g476B (.Q(g476B),.SE(test_seB),.SI(g440B),.D(g11338B),.CK(CKB));
SDFF_X1 U_g119B (.Q(g119B),.SE(test_seB),.SI(g476B),.D(g5918B),.CK(CKB));
SDFF_X1 U_g668B (.Q(g668B),.SE(test_seB),.SI(g119B),.D(g8922B),.CK(CKB));
SDFF_X1 U_g139B (.Q(g139B),.SE(test_seB),.SI(g668B),.D(g8049B),.CK(CKB));
SDFF_X1 U_g1149B (.Q(g1149B),.SE(test_seB),.SI(g139B),.D(g4342B),.CK(CKB));
SDFF_X1 U_g34B (.Q(g34B),.SE(test_seB),.SI(g1149B),.D(g10720B),.CK(CKB));
SDFF_X1 U_g1848B (.Q(g1848B),.SE(test_seB),.SI(g34B),.D(g6755B),.CK(CKB));
SDFF_X1 U_g263B (.Q(g263B),.SE(test_seB),.SI(g1848B),.D(g6897B),.CK(CKB));
SDFF_X1 U_g818B (.Q(g818B),.SE(test_seB),.SI(g263B),.D(g7709B),.CK(CKB));
SDFF_X1 U_g1747B (.Q(g1747B),.SE(test_seB),.SI(g818B),.D(g4255B),.CK(CKB));
SDFF_X1 U_g802B (.Q(g802B),.SE(test_seB),.SI(g1747B),.D(g5543B),.CK(CKB));
SDFF_X1 U_g275B (.Q(g275B),.SE(test_seB),.SI(g802B),.D(g6915B),.CK(CKB));
SDFF_X1 U_g1524B (.Q(g1524B),.SE(test_seB),.SI(g275B),.D(g6513B),.CK(CKB));
SDFF_X1 U_g1577B (.Q(g1577B),.SE(test_seB),.SI(g1524B),.D(g6480B),.CK(CKB));
SDFF_X1 U_g810B (.Q(g810B),.SE(test_seB),.SI(g1577B),.D(g6733B),.CK(CKB));
SDFF_X1 U_g391B (.Q(g391B),.SE(test_seB),.SI(g810B),.D(g11264B),.CK(CKB));
SDFF_X1 U_g658B (.Q(g658B),.SE(test_seB),.SI(g391B),.D(g8973B),.CK(CKB));
SDFF_X1 U_g1386B (.Q(g1386B),.SE(test_seB),.SI(g658B),.D(g6833B),.CK(CKB));
SDFF_X1 U_g253B (.Q(g253B),.SE(test_seB),.SI(g1386B),.D(g5996B),.CK(CKB));
SDFF_X1 U_g875B (.Q(g875B),.SE(test_seB),.SI(g253B),.D(g9508B),.CK(CKB));
SDFF_X1 U_g1125B (.Q(g1125B),.SE(test_seB),.SI(g875B),.D(g4473B),.CK(CKB));
SDFF_X1 U_g201B (.Q(g201B),.SE(test_seB),.SI(g1125B),.D(g5755B),.CK(CKB));
SDFF_X1 U_g1280B (.Q(g1280B),.SE(test_seB),.SI(g201B),.D(g7295B),.CK(CKB));
SDFF_X1 U_g1083B (.Q(g1083B),.SE(test_seB),.SI(g1280B),.D(g6068B),.CK(CKB));
SDFF_X1 U_g650B (.Q(g650B),.SE(test_seB),.SI(g1083B),.D(g7137B),.CK(CKB));
SDFF_X1 U_g1636B (.Q(g1636B),.SE(test_seB),.SI(g650B),.D(g8779B),.CK(CKB));
SDFF_X1 U_g853B (.Q(g853B),.SE(test_seB),.SI(g1636B),.D(g818B),.CK(CKB));
SDFF_X1 U_g421B (.Q(g421B),.SE(test_seB),.SI(g853B),.D(g11270B),.CK(CKB));
SDFF_X1 U_g762B (.Q(g762B),.SE(test_seB),.SI(g421B),.D(g5529B),.CK(CKB));
SDFF_X1 U_g956B (.Q(g956B),.SE(test_seB),.SI(g762B),.D(g11306B),.CK(CKB));
SDFF_X1 U_g378B (.Q(g378B),.SE(test_seB),.SI(g956B),.D(g11291B),.CK(CKB));
SDFF_X1 U_g1756B (.Q(g1756B),.SE(test_seB),.SI(g378B),.D(g4283B),.CK(CKB));
SDFF_X1 U_g589B (.Q(g589B),.SE(test_seB),.SI(g1756B),.D(g29B),.CK(CKB));
SDFF_X1 U_g841B (.Q(g841B),.SE(test_seB),.SI(g589B),.D(g806B),.CK(CKB));
SDFF_X1 U_g1027B (.Q(g1027B),.SE(test_seB),.SI(g841B),.D(g6894B),.CK(CKB));
SDFF_X1 U_g1003B (.Q(g1003B),.SE(test_seB),.SI(g1027B),.D(g6902B),.CK(CKB));
SDFF_X1 U_g1403B (.Q(g1403B),.SE(test_seB),.SI(g1003B),.D(g8765B),.CK(CKB));
SDFF_X1 U_g1145B (.Q(g1145B),.SE(test_seB),.SI(g1403B),.D(g4498B),.CK(CKB));
SDFF_X1 U_g1107B (.Q(g1107B),.SE(test_seB),.SI(g1145B),.D(g5148B),.CK(CKB));
SDFF_X1 U_g1223B (.Q(g1223B),.SE(test_seB),.SI(g1107B),.D(g7581B),.CK(CKB));
SDFF_X1 U_g406B (.Q(g406B),.SE(test_seB),.SI(g1223B),.D(g11267B),.CK(CKB));
SDFF_X1 U_g1811B (.Q(g1811B),.SE(test_seB),.SI(g406B),.D(g10936B),.CK(CKB));
SDFF_X1 U_g1642B (.Q(g1642B),.SE(test_seB),.SI(g1811B),.D(g10784B),.CK(CKB));
SDFF_X1 U_g1047B (.Q(g1047B),.SE(test_seB),.SI(g1642B),.D(g7211B),.CK(CKB));
SDFF_X1 U_g1654B (.Q(g1654B),.SE(test_seB),.SI(g1047B),.D(g10765B),.CK(CKB));
SDFF_X1 U_g197B (.Q(g197B),.SE(test_seB),.SI(g1654B),.D(g6332B),.CK(CKB));
SDFF_X1 U_g1595B (.Q(g1595B),.SE(test_seB),.SI(g197B),.D(g6479B),.CK(CKB));
SDFF_X1 U_g1537B (.Q(g1537B),.SE(test_seB),.SI(g1595B),.D(g6537B),.CK(CKB));
SDFF_X1 U_g727B (.Q(g727B),.SE(test_seB),.SI(g1537B),.D(g8434B),.CK(CKB));
SDFF_X1 U_g999B (.Q(g999B),.SE(test_seB),.SI(g727B),.D(g6908B),.CK(CKB));
SDFF_X1 U_g798B (.Q(g798B),.SE(test_seB),.SI(g999B),.D(g6243B),.CK(CKB));
SDFF_X1 U_g481B (.Q(g481B),.SE(test_seB),.SI(g798B),.D(g11324B),.CK(CKB));
SDFF_X1 U_g754B (.Q(g754B),.SE(test_seB),.SI(g481B),.D(g3462B),.CK(CKB));
SDFF_X1 U_g1330B (.Q(g1330B),.SE(test_seB),.SI(g754B),.D(g11609B),.CK(CKB));
SDFF_X1 U_g845B (.Q(g845B),.SE(test_seB),.SI(g1330B),.D(g810B),.CK(CKB));
SDFF_X1 U_g790B (.Q(g790B),.SE(test_seB),.SI(g845B),.D(g8244B),.CK(CKB));
SDFF_X1 U_g1512B (.Q(g1512B),.SE(test_seB),.SI(g790B),.D(g8194B),.CK(CKB));
SDFF_X1 U_g114B (.Q(g114B),.SE(test_seB),.SI(g1512B),.D(g113B),.CK(CKB));
SDFF_X1 U_g1490B (.Q(g1490B),.SE(test_seB),.SI(g114B),.D(g8052B),.CK(CKB));
SDFF_X1 U_g1166B (.Q(g1166B),.SE(test_seB),.SI(g1490B),.D(g4325B),.CK(CKB));
SDFF_X1 U_g1056B (.Q(g1056B),.SE(test_seB),.SI(g1166B),.D(g7231B),.CK(CKB));
SDFF_X1 U_g348B (.Q(g348B),.SE(test_seB),.SI(g1056B),.D(g11481B),.CK(CKB));
SDFF_X1 U_g868B (.Q(g868B),.SE(test_seB),.SI(g348B),.D(g874B),.CK(CKB));
SDFF_X1 U_g1260B (.Q(g1260B),.SE(test_seB),.SI(g868B),.D(g7301B),.CK(CKB));
SDFF_X1 U_g260B (.Q(g260B),.SE(test_seB),.SI(g1260B),.D(g6035B),.CK(CKB));
SDFF_X1 U_g131B (.Q(g131B),.SE(test_seB),.SI(g260B),.D(g8059B),.CK(CKB));
SDFF_X1 U_g7B (.Q(g7B),.SE(test_seB),.SI(g131B),.D(g1854B),.CK(CKB));
SDFF_X1 U_g258B (.Q(g258B),.SE(test_seB),.SI(g7B),.D(g6015B),.CK(CKB));
SDFF_X1 U_g521B (.Q(g521B),.SE(test_seB),.SI(g258B),.D(g11330B),.CK(CKB));
SDFF_X1 U_g1318B (.Q(g1318B),.SE(test_seB),.SI(g521B),.D(g11605B),.CK(CKB));
SDFF_X1 U_g1872B (.Q(g1872B),.SE(test_seB),.SI(g1318B),.D(g8921B),.CK(CKB));
SDFF_X1 U_g677B (.Q(g677B),.SE(test_seB),.SI(g1872B),.D(g8883B),.CK(CKB));
SDFF_X1 U_g582B (.Q(g582B),.SE(test_seB),.SI(g677B),.D(g28B),.CK(CKB));
SDFF_X1 U_g1393B (.Q(g1393B),.SE(test_seB),.SI(g582B),.D(g6163B),.CK(CKB));
SDFF_X1 U_g1549B (.Q(g1549B),.SE(test_seB),.SI(g1393B),.D(g6523B),.CK(CKB));
SDFF_X1 U_g947B (.Q(g947B),.SE(test_seB),.SI(g1549B),.D(g11300B),.CK(CKB));
SDFF_X1 U_g1834B (.Q(g1834B),.SE(test_seB),.SI(g947B),.D(g9555B),.CK(CKB));
SDFF_X1 U_g1598B (.Q(g1598B),.SE(test_seB),.SI(g1834B),.D(g6481B),.CK(CKB));
SDFF_X1 U_g1121B (.Q(g1121B),.SE(test_seB),.SI(g1598B),.D(g4471B),.CK(CKB));
SDFF_X1 U_g1321B (.Q(g1321B),.SE(test_seB),.SI(g1121B),.D(g11606B),.CK(CKB));
SDFF_X1 U_g506B (.Q(g506B),.SE(test_seB),.SI(g1321B),.D(g11335B),.CK(CKB));
SDFF_X1 U_g546B (.Q(g546B),.SE(test_seB),.SI(g506B),.D(g10791B),.CK(CKB));
SDFF_X1 U_g1909B (.Q(g1909B),.SE(test_seB),.SI(g546B),.D(g8939B),.CK(CKB));
SDFF_X1 U_g755B (.Q(g755B),.SE(test_seB),.SI(g1909B),.D(g83B),.CK(CKB));
SDFF_X1 U_g1552B (.Q(g1552B),.SE(test_seB),.SI(g755B),.D(g6529B),.CK(CKB));
SDFF_X1 U_g584B (.Q(g584B),.SE(test_seB),.SI(g1552B),.D(g101B),.CK(CKB));
SDFF_X1 U_g1687B (.Q(g1687B),.SE(test_seB),.SI(g584B),.D(g10776B),.CK(CKB));
SDFF_X1 U_g1586B (.Q(g1586B),.SE(test_seB),.SI(g1687B),.D(g6514B),.CK(CKB));
SDFF_X1 U_g324B (.Q(g324B),.SE(test_seB),.SI(g1586B),.D(g259B),.CK(CKB));
SDFF_X1 U_g1141B (.Q(g1141B),.SE(test_seB),.SI(g324B),.D(g4490B),.CK(CKB));
SDFF_X1 U_g1570B (.Q(g1570B),.SE(test_seB),.SI(g1141B),.D(I8503B),.CK(CKB));
SDFF_X1 U_g1341B (.Q(g1341B),.SE(test_seB),.SI(g1570B),.D(g11639B),.CK(CKB));
SDFF_X1 U_g1710B (.Q(g1710B),.SE(test_seB),.SI(g1341B),.D(g4089B),.CK(CKB));
SDFF_X1 U_g1645B (.Q(g1645B),.SE(test_seB),.SI(g1710B),.D(g10785B),.CK(CKB));
SDFF_X1 U_g115B (.Q(g115B),.SE(test_seB),.SI(g1645B),.D(g6179B),.CK(CKB));
SDFF_X1 U_g135B (.Q(g135B),.SE(test_seB),.SI(g115B),.D(g8053B),.CK(CKB));
SDFF_X1 U_g525B (.Q(g525B),.SE(test_seB),.SI(g135B),.D(g11329B),.CK(CKB));
SDFF_X1 U_g581B (.Q(g581B),.SE(test_seB),.SI(g525B),.D(g104B),.CK(CKB));
SDFF_X1 U_g1607B (.Q(g1607B),.SE(test_seB),.SI(g581B),.D(g6515B),.CK(CKB));
SDFF_X1 U_g321B (.Q(g321B),.SE(test_seB),.SI(g1607B),.D(g258B),.CK(CKB));
SDFF_X1 U_g67B (.Q(g67B),.SE(test_seB),.SI(g321B),.D(g7204B),.CK(CKB));
SDFF_X1 U_g1275B (.Q(g1275B),.SE(test_seB),.SI(g67B),.D(g11443B),.CK(CKB));
SDFF_X1 U_g1311B (.Q(g1311B),.SE(test_seB),.SI(g1275B),.D(g11603B),.CK(CKB));
SDFF_X1 U_g1615B (.Q(g1615B),.SE(test_seB),.SI(g1311B),.D(g8770B),.CK(CKB));
SDFF_X1 U_g382B (.Q(g382B),.SE(test_seB),.SI(g1615B),.D(g11292B),.CK(CKB));
SDFF_X1 U_g1374B (.Q(g1374B),.SE(test_seB),.SI(g382B),.D(g6331B),.CK(CKB));
SDFF_X1 U_g266B (.Q(g266B),.SE(test_seB),.SI(g1374B),.D(g6900B),.CK(CKB));
SDFF_X1 U_g1284B (.Q(g1284B),.SE(test_seB),.SI(g266B),.D(g7294B),.CK(CKB));
SDFF_X1 U_g1380B (.Q(g1380B),.SE(test_seB),.SI(g1284B),.D(g6829B),.CK(CKB));
SDFF_X1 U_g673B (.Q(g673B),.SE(test_seB),.SI(g1380B),.D(g8428B),.CK(CKB));
SDFF_X1 U_g1853B (.Q(g1853B),.SE(test_seB),.SI(g673B),.D(g4904B),.CK(CKB));
SDFF_X1 U_g162B (.Q(g162B),.SE(test_seB),.SI(g1853B),.D(g8054B),.CK(CKB));
SDFF_X1 U_g411B (.Q(g411B),.SE(test_seB),.SI(g162B),.D(g11268B),.CK(CKB));
SDFF_X1 U_g431B (.Q(g431B),.SE(test_seB),.SI(g411B),.D(g11262B),.CK(CKB));
SDFF_X1 U_g1905B (.Q(g1905B),.SE(test_seB),.SI(g431B),.D(g8283B),.CK(CKB));
SDFF_X1 U_g1515B (.Q(g1515B),.SE(test_seB),.SI(g1905B),.D(g6193B),.CK(CKB));
SDFF_X1 U_g1630B (.Q(g1630B),.SE(test_seB),.SI(g1515B),.D(g8776B),.CK(CKB));
SDFF_X1 U_g49B (.Q(g49B),.SE(test_seB),.SI(g1630B),.D(g7143B),.CK(CKB));
SDFF_X1 U_g991B (.Q(g991B),.SE(test_seB),.SI(g49B),.D(g6898B),.CK(CKB));
SDFF_X1 U_g1300B (.Q(g1300B),.SE(test_seB),.SI(g991B),.D(g7291B),.CK(CKB));
SDFF_X1 U_g339B (.Q(g339B),.SE(test_seB),.SI(g1300B),.D(g11478B),.CK(CKB));
SDFF_X1 U_g256B (.Q(g256B),.SE(test_seB),.SI(g339B),.D(g6000B),.CK(CKB));
SDFF_X1 U_g1750B (.Q(g1750B),.SE(test_seB),.SI(g256B),.D(g4264B),.CK(CKB));
SDFF_X1 U_g585B (.Q(g585B),.SE(test_seB),.SI(g1750B),.D(g102B),.CK(CKB));
SDFF_X1 U_g1440B (.Q(g1440B),.SE(test_seB),.SI(g585B),.D(g8768B),.CK(CKB));
SDFF_X1 U_g1666B (.Q(g1666B),.SE(test_seB),.SI(g1440B),.D(g10863B),.CK(CKB));
SDFF_X1 U_g1528B (.Q(g1528B),.SE(test_seB),.SI(g1666B),.D(g6522B),.CK(CKB));
SDFF_X1 U_g1351B (.Q(g1351B),.SE(test_seB),.SI(g1528B),.D(g11641B),.CK(CKB));
SDFF_X1 U_g1648B (.Q(g1648B),.SE(test_seB),.SI(g1351B),.D(g10780B),.CK(CKB));
SDFF_X1 U_g127B (.Q(g127B),.SE(test_seB),.SI(g1648B),.D(g8044B),.CK(CKB));
SDFF_X1 U_g1618B (.Q(g1618B),.SE(test_seB),.SI(g127B),.D(g11579B),.CK(CKB));
SDFF_X1 U_g1235B (.Q(g1235B),.SE(test_seB),.SI(g1618B),.D(g7296B),.CK(CKB));
SDFF_X1 U_g299B (.Q(g299B),.SE(test_seB),.SI(g1235B),.D(g6923B),.CK(CKB));
SDFF_X1 U_g435B (.Q(g435B),.SE(test_seB),.SI(g299B),.D(g11261B),.CK(CKB));
SDFF_X1 U_g64B (.Q(g64B),.SE(test_seB),.SI(g435B),.D(g6638B),.CK(CKB));
SDFF_X1 U_g1555B (.Q(g1555B),.SE(test_seB),.SI(g64B),.D(g6534B),.CK(CKB));
SDFF_X1 U_g995B (.Q(g995B),.SE(test_seB),.SI(g1555B),.D(g6895B),.CK(CKB));
SDFF_X1 U_g1621B (.Q(g1621B),.SE(test_seB),.SI(g995B),.D(g8771B),.CK(CKB));
SDFF_X1 U_g1113B (.Q(g1113B),.SE(test_seB),.SI(g1621B),.D(g4506B),.CK(CKB));
SDFF_X1 U_g643B (.Q(g643B),.SE(test_seB),.SI(g1113B),.D(g7441B),.CK(CKB));
SDFF_X1 U_g1494B (.Q(g1494B),.SE(test_seB),.SI(g643B),.D(g8055B),.CK(CKB));
SDFF_X1 U_g1567B (.Q(g1567B),.SE(test_seB),.SI(g1494B),.D(g6468B),.CK(CKB));
SDFF_X1 U_g691B (.Q(g691B),.SE(test_seB),.SI(g1567B),.D(g8430B),.CK(CKB));
SDFF_X1 U_g534B (.Q(g534B),.SE(test_seB),.SI(g691B),.D(g11327B),.CK(CKB));
SDFF_X1 U_g1776B (.Q(g1776B),.SE(test_seB),.SI(g534B),.D(g6508B),.CK(CKB));
SDFF_X1 U_g569B (.Q(g569B),.SE(test_seB),.SI(g1776B),.D(g10717B),.CK(CKB));
SDFF_X1 U_g1160B (.Q(g1160B),.SE(test_seB),.SI(g569B),.D(g4334B),.CK(CKB));
SDFF_X1 U_g1360B (.Q(g1360B),.SE(test_seB),.SI(g1160B),.D(g9526B),.CK(CKB));
SDFF_X1 U_g1050B (.Q(g1050B),.SE(test_seB),.SI(g1360B),.D(g7218B),.CK(CKB));
SDFF_X1 U_g1B (.Q(g1B),.SE(test_seB),.SI(g1050B),.D(g6679B),.CK(CKB));
SDFF_X1 U_g511B (.Q(g511B),.SE(test_seB),.SI(g1B),.D(g11336B),.CK(CKB));
SDFF_X1 U_g1724B (.Q(g1724B),.SE(test_seB),.SI(g511B),.D(g10771B),.CK(CKB));
SDFF_X1 U_g12B (.Q(g12B),.SE(test_seB),.SI(g1724B),.D(g5445B),.CK(CKB));
SDFF_X1 U_g1878B (.Q(g1878B),.SE(test_seB),.SI(g12B),.D(g8559B),.CK(CKB));
SDFF_X1 U_g73B (.Q(g73B),.SE(test_seB),.SI(g1878B),.D(g7219B),.CK(CKB));
INV_X1 FE_OFC370_g4525C (.ZN(FE_OFN370_g4525C),.A(FE_OFN368_g4525C));
INV_X1 FE_OFC369_g4525C (.ZN(FE_OFN369_g4525C),.A(FE_OFN368_g4525C));
INV_X1 FE_OFC368_g4525C (.ZN(FE_OFN368_g4525C),.A(FE_OFN362_g4525C));
BUF_X3 FE_OFC367_g3521C (.Z(FE_OFN367_g3521C),.A(FE_OFN366_g3521C));
BUF_X3 FE_OFC366_g3521C (.Z(FE_OFN366_g3521C),.A(FE_OFN358_g3521C));
BUF_X3 FE_OFC365_g5361C (.Z(FE_OFN365_g5361C),.A(FE_OFN356_g5361C));
BUF_X3 FE_OFC364_g3015C (.Z(FE_OFN364_g3015C),.A(FE_OFN348_g3015C));
BUF_X3 FE_OFC363_I5565C (.Z(FE_OFN363_I5565C),.A(FE_OFN343_I5565C));
INV_X1 FE_OFC362_g4525C (.ZN(FE_OFN362_g4525C),.A(FE_OFN360_g4525C));
INV_X1 FE_OFC360_g4525C (.ZN(FE_OFN360_g4525C),.A(FE_OFN339_g4525C));
BUF_X3 FE_OFC359_g18C (.Z(FE_OFN359_g18C),.A(FE_OFN324_g18C));
BUF_X3 FE_OFC358_g3521C (.Z(FE_OFN358_g3521C),.A(g3521C));
BUF_X3 FE_OFC357_g3521C (.Z(FE_OFN357_g3521C),.A(FE_OFN366_g3521C));
INV_X1 FE_OFC356_g5361C (.ZN(FE_OFN356_g5361C),.A(FE_OFN354_g5361C));
INV_X1 FE_OFC354_g5361C (.ZN(FE_OFN354_g5361C),.A(FE_OFN318_g5361C));
BUF_X3 FE_OFC353_g5117C (.Z(FE_OFN353_g5117C),.A(FE_OFN315_g5117C));
BUF_X3 FE_OFC352_g109C (.Z(FE_OFN352_g109C),.A(FE_OFN269_g109C));
BUF_X3 FE_OFC351_g3913C (.Z(FE_OFN351_g3913C),.A(FE_OFN302_g3913C));
BUF_X3 FE_OFC350_g3121C (.Z(FE_OFN350_g3121C),.A(FE_OFN155_g3121C));
BUF_X3 FE_OFC349_I6424C (.Z(FE_OFN349_I6424C),.A(FE_OFN308_I6424C));
BUF_X3 FE_OFC348_g3015C (.Z(FE_OFN348_g3015C),.A(FE_OFN298_g3015C));
BUF_X3 FE_OFC347_g3914C (.Z(FE_OFN347_g3914C),.A(FE_OFN296_g3914C));
BUF_X3 FE_OFC346_g4381C (.Z(FE_OFN346_g4381C),.A(g4381C));
BUF_X3 FE_OFC345_g3015C (.Z(FE_OFN345_g3015C),.A(FE_OFN297_g3015C));
BUF_X3 FE_OFC344_g3586C (.Z(FE_OFN344_g3586C),.A(FE_OFN287_g3586C));
INV_X1 FE_OFC343_I5565C (.ZN(FE_OFN343_I5565C),.A(FE_OFN340_I5565C));
INV_X1 FE_OFC340_I5565C (.ZN(FE_OFN340_I5565C),.A(FE_OFN233_I5565C));
INV_X1 FE_OFC339_g4525C (.ZN(FE_OFN339_g4525C),.A(FE_OFN337_g4525C));
INV_X1 FE_OFC337_g4525C (.ZN(FE_OFN337_g4525C),.A(g4525C));
BUF_X3 FE_OFC336_g1690C (.Z(FE_OFN336_g1690C),.A(FE_OFN245_g1690C));
BUF_X3 FE_OFC335_g4737C (.Z(FE_OFN335_g4737C),.A(g4737C));
BUF_X3 FE_OFC334_g7045C (.Z(FE_OFN334_g7045C),.A(g7045C));
BUF_X3 FE_OFC333_g4294C (.Z(FE_OFN333_g4294C),.A(g4294C));
BUF_X3 FE_OFC332_g8748C (.Z(FE_OFN332_g8748C),.A(g8748C));
BUF_X3 FE_OFC331_g8696C (.Z(FE_OFN331_g8696C),.A(g8696C));
BUF_X3 FE_OFC330_g7638C (.Z(FE_OFN330_g7638C),.A(FE_OFN189_g7638C));
BUF_X3 FE_OFC329_g8763C (.Z(FE_OFN329_g8763C),.A(g8763C));
BUF_X3 FE_OFC328_g8709C (.Z(FE_OFN328_g8709C),.A(g8709C));
BUF_X3 FE_OFC325_g18C (.Z(FE_OFN325_g18C),.A(FE_OFN359_g18C));
BUF_X3 FE_OFC324_g18C (.Z(FE_OFN324_g18C),.A(FE_OFN260_g18C));
BUF_X3 FE_OFC322_g4449C (.Z(FE_OFN322_g4449C),.A(g4449C));
BUF_X3 FE_OFC321_g5261C (.Z(FE_OFN321_g5261C),.A(g5261C));
BUF_X3 FE_OFC320_g5361C (.Z(FE_OFN320_g5361C),.A(FE_OFN319_g5361C));
BUF_X3 FE_OFC319_g5361C (.Z(FE_OFN319_g5361C),.A(FE_OFN166_g5361C));
INV_X1 FE_OFC318_g5361C (.ZN(FE_OFN318_g5361C),.A(FE_OFN316_g5361C));
INV_X1 FE_OFC316_g5361C (.ZN(FE_OFN316_g5361C),.A(FE_OFN168_g5361C));
INV_X1 FE_OFC315_g5117C (.ZN(FE_OFN315_g5117C),.A(FE_OFN312_g5117C));
INV_X1 FE_OFC312_g5117C (.ZN(FE_OFN312_g5117C),.A(g5117C));
BUF_X3 FE_OFC310_g4336C (.Z(FE_OFN310_g4336C),.A(g4336C));
BUF_X3 FE_OFC308_I6424C (.Z(FE_OFN308_I6424C),.A(FE_OFN160_I6424C));
BUF_X3 FE_OFC307_g4010C (.Z(FE_OFN307_g4010C),.A(g4010C));
BUF_X3 FE_OFC306_g5128C (.Z(FE_OFN306_g5128C),.A(g5128C));
BUF_X3 FE_OFC305_g5151C (.Z(FE_OFN305_g5151C),.A(FE_OFN304_g5151C));
BUF_X3 FE_OFC304_g5151C (.Z(FE_OFN304_g5151C),.A(FE_OFN176_g5151C));
BUF_X3 FE_OFC303_g4678C (.Z(FE_OFN303_g4678C),.A(g4678C));
BUF_X3 FE_OFC302_g3913C (.Z(FE_OFN302_g3913C),.A(g3913C));
BUF_X3 FE_OFC300_g4002C (.Z(FE_OFN300_g4002C),.A(g4002C));
BUF_X3 FE_OFC299_g4457C (.Z(FE_OFN299_g4457C),.A(g4457C));
BUF_X3 FE_OFC298_g3015C (.Z(FE_OFN298_g3015C),.A(FE_OFN119_g3015C));
BUF_X3 FE_OFC297_g3015C (.Z(FE_OFN297_g3015C),.A(FE_OFN348_g3015C));
INV_X1 FE_OFC296_g3914C (.ZN(FE_OFN296_g3914C),.A(FE_OFN294_g3914C));
INV_X1 FE_OFC294_g3914C (.ZN(FE_OFN294_g3914C),.A(FE_OFN113_g3914C));
BUF_X3 FE_OFC293_g3015C (.Z(FE_OFN293_g3015C),.A(FE_OFN292_g3015C));
BUF_X3 FE_OFC292_g3015C (.Z(FE_OFN292_g3015C),.A(FE_OFN345_g3015C));
BUF_X3 FE_OFC291_g4880C (.Z(FE_OFN291_g4880C),.A(FE_OFN290_g4880C));
BUF_X3 FE_OFC290_g4880C (.Z(FE_OFN290_g4880C),.A(g4880C));
BUF_X3 FE_OFC289_g4679C (.Z(FE_OFN289_g4679C),.A(g4679C));
BUF_X3 FE_OFC288_g4263C (.Z(FE_OFN288_g4263C),.A(g4263C));
INV_X1 FE_OFC287_g3586C (.ZN(FE_OFN287_g3586C),.A(FE_OFN284_g3586C));
INV_X1 FE_OFC284_g3586C (.ZN(FE_OFN284_g3586C),.A(FE_OFN110_g3586C));
BUF_X3 FE_OFC283_I8869C (.Z(FE_OFN283_I8869C),.A(FE_OFN97_I8869C));
BUF_X3 FE_OFC282_g6165C (.Z(FE_OFN282_g6165C),.A(g6165C));
BUF_X3 FE_OFC281_g2216C (.Z(FE_OFN281_g2216C),.A(FE_OFN95_g2216C));
BUF_X3 FE_OFC280_g9536C (.Z(FE_OFN280_g9536C),.A(FE_OFN64_g9536C));
BUF_X3 FE_OFC279_g11157C (.Z(FE_OFN279_g11157C),.A(g11157C));
BUF_X3 FE_OFC278_g10927C (.Z(FE_OFN278_g10927C),.A(g10927C));
BUF_X3 FE_OFC277_g48C (.Z(FE_OFN277_g48C),.A(FE_OFN276_g48C));
BUF_X3 FE_OFC276_g48C (.Z(FE_OFN276_g48C),.A(FE_OFN275_g48C));
BUF_X3 FE_OFC275_g48C (.Z(FE_OFN275_g48C),.A(g48C));
BUF_X3 FE_OFC273_g85C (.Z(FE_OFN273_g85C),.A(FE_OFN271_g85C));
BUF_X3 FE_OFC271_g85C (.Z(FE_OFN271_g85C),.A(g85C));
BUF_X3 FE_OFC269_g109C (.Z(FE_OFN269_g109C),.A(FE_OFN267_g109C));
BUF_X3 FE_OFC267_g109C (.Z(FE_OFN267_g109C),.A(g109C));
BUF_X3 FE_OFC266_g18C (.Z(FE_OFN266_g18C),.A(FE_OFN325_g18C));
BUF_X3 FE_OFC260_g18C (.Z(FE_OFN260_g18C),.A(g2355C));
BUF_X3 FE_OFC254_g461C (.Z(FE_OFN254_g461C),.A(g461C));
BUF_X3 FE_OFC253_g1786C (.Z(FE_OFN253_g1786C),.A(g1786C));
BUF_X3 FE_OFC252_g1791C (.Z(FE_OFN252_g1791C),.A(g1791C));
BUF_X3 FE_OFC251_g1801C (.Z(FE_OFN251_g1801C),.A(g1801C));
BUF_X3 FE_OFC250_g471C (.Z(FE_OFN250_g471C),.A(g471C));
BUF_X3 FE_OFC248_g466C (.Z(FE_OFN248_g466C),.A(g466C));
BUF_X3 FE_OFC247_g1771C (.Z(FE_OFN247_g1771C),.A(g1771C));
INV_X1 FE_OFC245_g1690C (.ZN(FE_OFN245_g1690C),.A(g2424C));
BUF_X3 FE_OFC241_g1690C (.Z(FE_OFN241_g1690C),.A(g1690C));
BUF_X3 FE_OFC240_g1110C (.Z(FE_OFN240_g1110C),.A(g1110C));
BUF_X3 FE_OFC239_g1796C (.Z(FE_OFN239_g1796C),.A(g1796C));
BUF_X3 FE_OFC238_g1781C (.Z(FE_OFN238_g1781C),.A(g1781C));
BUF_X3 FE_OFC237_g1806C (.Z(FE_OFN237_g1806C),.A(g1806C));
BUF_X3 FE_OFC236_g1776C (.Z(FE_OFN236_g1776C),.A(g1776C));
BUF_X3 FE_OFC235_g2024C (.Z(FE_OFN235_g2024C),.A(FE_OFN234_g2024C));
BUF_X3 FE_OFC234_g2024C (.Z(FE_OFN234_g2024C),.A(g2024C));
INV_X1 FE_OFC233_I5565C (.ZN(FE_OFN233_I5565C),.A(FE_OFN230_I5565C));
INV_X1 FE_OFC230_I5565C (.ZN(FE_OFN230_I5565C),.A(I6360C));
INV_X1 FE_OFC229_g3880C (.ZN(FE_OFN229_g3880C),.A(FE_OFN227_g3880C));
INV_X1 FE_OFC227_g3880C (.ZN(FE_OFN227_g3880C),.A(FE_OFN226_g3880C));
BUF_X3 FE_OFC226_g3880C (.Z(FE_OFN226_g3880C),.A(g3880C));
BUF_X3 FE_OFC225_g2276C (.Z(FE_OFN225_g2276C),.A(FE_OFN224_g2276C));
BUF_X3 FE_OFC224_g2276C (.Z(FE_OFN224_g2276C),.A(g2276C));
BUF_X3 FE_OFC223_g4401C (.Z(FE_OFN223_g4401C),.A(g4401C));
BUF_X3 FE_OFC221_g3440C (.Z(FE_OFN221_g3440C),.A(g3440C));
BUF_X3 FE_OFC219_g5557C (.Z(FE_OFN219_g5557C),.A(FE_OFN218_g5557C));
BUF_X3 FE_OFC218_g5557C (.Z(FE_OFN218_g5557C),.A(g5557C));
INV_X1 FE_OFC217_g5013C (.ZN(FE_OFN217_g5013C),.A(g6403C));
BUF_X3 FE_OFC213_g6003C (.Z(FE_OFN213_g6003C),.A(g6003C));
BUF_X3 FE_OFC211_g7246C (.Z(FE_OFN211_g7246C),.A(FE_OFN210_g7246C));
BUF_X3 FE_OFC210_g7246C (.Z(FE_OFN210_g7246C),.A(g7246C));
INV_X1 FE_OFC209_g6863C (.ZN(FE_OFN209_g6863C),.A(FE_OFN207_g6863C));
INV_X1 FE_OFC207_g6863C (.ZN(FE_OFN207_g6863C),.A(FE_OFN206_g6863C));
BUF_X3 FE_OFC206_g6863C (.Z(FE_OFN206_g6863C),.A(g6863C));
BUF_X3 FE_OFC204_g3664C (.Z(FE_OFN204_g3664C),.A(g3664C));
BUF_X3 FE_OFC200_g4921C (.Z(FE_OFN200_g4921C),.A(g4921C));
BUF_X3 FE_OFC199_g7697C (.Z(FE_OFN199_g7697C),.A(FE_OFN198_g7697C));
INV_X1 FE_OFC198_g7697C (.ZN(FE_OFN198_g7697C),.A(FE_OFN196_g7697C));
INV_X1 FE_OFC196_g7697C (.ZN(FE_OFN196_g7697C),.A(g7697C));
INV_X1 FE_OFC195_g6488C (.ZN(FE_OFN195_g6488C),.A(FE_OFN192_g6488C));
INV_X1 FE_OFC192_g6488C (.ZN(FE_OFN192_g6488C),.A(g6488C));
BUF_X3 FE_OFC191_g6488C (.Z(FE_OFN191_g6488C),.A(g6488C));
INV_X1 FE_OFC189_g7638C (.ZN(FE_OFN189_g7638C),.A(FE_OFN187_g7638C));
INV_X1 FE_OFC187_g7638C (.ZN(FE_OFN187_g7638C),.A(g7638C));
BUF_X3 FE_OFC184_I7048C (.Z(FE_OFN184_I7048C),.A(I7048C));
BUF_X3 FE_OFC180_g5354C (.Z(FE_OFN180_g5354C),.A(FE_OFN179_g5354C));
BUF_X3 FE_OFC179_g5354C (.Z(FE_OFN179_g5354C),.A(FE_OFN178_g5354C));
BUF_X3 FE_OFC178_g5354C (.Z(FE_OFN178_g5354C),.A(g5354C));
BUF_X3 FE_OFC177_g5919C (.Z(FE_OFN177_g5919C),.A(g5919C));
BUF_X3 FE_OFC176_g5151C (.Z(FE_OFN176_g5151C),.A(FE_OFN306_g5128C));
INV_X1 FE_OFC168_g5361C (.ZN(FE_OFN168_g5361C),.A(FE_OFN166_g5361C));
INV_X1 FE_OFC166_g5361C (.ZN(FE_OFN166_g5361C),.A(FE_OFN164_g5361C));
INV_X1 FE_OFC164_g5361C (.ZN(FE_OFN164_g5361C),.A(FE_OFN161_g5361C));
INV_X1 FE_OFC161_g5361C (.ZN(FE_OFN161_g5361C),.A(g5361C));
BUF_X3 FE_OFC160_I6424C (.Z(FE_OFN160_I6424C),.A(FE_OFN350_g3121C));
BUF_X3 FE_OFC155_g3121C (.Z(FE_OFN155_g3121C),.A(g3121C));
BUF_X3 FE_OFC154_g4640C (.Z(FE_OFN154_g4640C),.A(FE_OFN153_g4640C));
INV_X1 FE_OFC153_g4640C (.ZN(FE_OFN153_g4640C),.A(FE_OFN321_g5261C));
BUF_X4 FE_OFC147_g4682C (.Z(FE_OFN147_g4682C),.A(FE_OFN146_g4682C));
BUF_X3 FE_OFC146_g4682C (.Z(FE_OFN146_g4682C),.A(FE_OFN144_g4682C));
INV_X1 FE_OFC144_g4682C (.ZN(FE_OFN144_g4682C),.A(FE_OFN142_g4682C));
INV_X1 FE_OFC142_g4682C (.ZN(FE_OFN142_g4682C),.A(g4682C));
INV_X1 FE_OFC141_g3829C (.ZN(FE_OFN141_g3829C),.A(FE_OFN299_g4457C));
BUF_X3 FE_OFC137_g3829C (.Z(FE_OFN137_g3829C),.A(g3829C));
INV_X1 FE_OFC136_g3863C (.ZN(FE_OFN136_g3863C),.A(FE_OFN134_g3863C));
INV_X1 FE_OFC134_g3863C (.ZN(FE_OFN134_g3863C),.A(g3863C));
BUF_X3 FE_OFC133_g3015C (.Z(FE_OFN133_g3015C),.A(FE_OFN131_g3015C));
BUF_X3 FE_OFC132_g3015C (.Z(FE_OFN132_g3015C),.A(FE_OFN293_g3015C));
INV_X1 FE_OFC131_g3015C (.ZN(FE_OFN131_g3015C),.A(FE_OFN291_g4880C));
BUF_X3 FE_OFC119_g3015C (.Z(FE_OFN119_g3015C),.A(g3015C));
BUF_X3 FE_OFC118_g4807C (.Z(FE_OFN118_g4807C),.A(FE_OFN117_g4807C));
BUF_X3 FE_OFC117_g4807C (.Z(FE_OFN117_g4807C),.A(FE_OFN116_g4807C));
BUF_X3 FE_OFC116_g4807C (.Z(FE_OFN116_g4807C),.A(FE_OFN115_g4807C));
BUF_X3 FE_OFC115_g4807C (.Z(FE_OFN115_g4807C),.A(g4807C));
INV_X1 FE_OFC113_g3914C (.ZN(FE_OFN113_g3914C),.A(FE_OFN111_g3914C));
INV_X1 FE_OFC111_g3914C (.ZN(FE_OFN111_g3914C),.A(g4673C));
INV_X1 FE_OFC110_g3586C (.ZN(FE_OFN110_g3586C),.A(g4263C));
BUF_X3 FE_OFC103_g3586C (.Z(FE_OFN103_g3586C),.A(FE_OFN102_g3586C));
BUF_X3 FE_OFC102_g3586C (.Z(FE_OFN102_g3586C),.A(g3586C));
BUF_X3 FE_OFC100_g4421C (.Z(FE_OFN100_g4421C),.A(FE_OFN99_g4421C));
BUF_X3 FE_OFC99_g4421C (.Z(FE_OFN99_g4421C),.A(g4421C));
BUF_X3 FE_OFC97_I8869C (.Z(FE_OFN97_I8869C),.A(I8869C));
BUF_X3 FE_OFC96_g2169C (.Z(FE_OFN96_g2169C),.A(g2169C));
BUF_X3 FE_OFC95_g2216C (.Z(FE_OFN95_g2216C),.A(FE_OFN93_g2216C));
BUF_X3 FE_OFC93_g2216C (.Z(FE_OFN93_g2216C),.A(FE_OFN92_g2216C));
BUF_X3 FE_OFC92_g2216C (.Z(FE_OFN92_g2216C),.A(g2216C));
BUF_X3 FE_OFC91_g2172C (.Z(FE_OFN91_g2172C),.A(g2172C));
BUF_X3 FE_OFC90_I11360C (.Z(FE_OFN90_I11360C),.A(FE_OFN89_I11360C));
BUF_X3 FE_OFC89_I11360C (.Z(FE_OFN89_I11360C),.A(I11360C));
BUF_X3 FE_OFC88_g2178C (.Z(FE_OFN88_g2178C),.A(g2178C));
BUF_X3 FE_OFC87_g2176C (.Z(FE_OFN87_g2176C),.A(FE_OFN86_g2176C));
BUF_X3 FE_OFC86_g2176C (.Z(FE_OFN86_g2176C),.A(FE_OFN85_g2176C));
BUF_X3 FE_OFC85_g2176C (.Z(FE_OFN85_g2176C),.A(FE_OFN83_g2176C));
INV_X1 FE_OFC84_g2176C (.ZN(FE_OFN84_g2176C),.A(FE_OFN81_g2176C));
INV_X1 FE_OFC83_g2176C (.ZN(FE_OFN83_g2176C),.A(FE_OFN81_g2176C));
INV_X1 FE_OFC82_g2176C (.ZN(FE_OFN82_g2176C),.A(FE_OFN81_g2176C));
INV_X1 FE_OFC81_g2176C (.ZN(FE_OFN81_g2176C),.A(g2176C));
BUF_X3 FE_OFC80_g2175C (.Z(FE_OFN80_g2175C),.A(g2175C));
INV_X1 FE_OFC79_g8700C (.ZN(FE_OFN79_g8700C),.A(g9097C));
BUF_X3 FE_OFC76_g8700C (.Z(FE_OFN76_g8700C),.A(g8700C));
BUF_X3 FE_OFC73_g8858C (.Z(FE_OFN73_g8858C),.A(g8858C));
BUF_X3 FE_OFC72_g9292C (.Z(FE_OFN72_g9292C),.A(FE_OFN71_g9292C));
BUF_X3 FE_OFC71_g9292C (.Z(FE_OFN71_g9292C),.A(g9292C));
BUF_X3 FE_OFC70_g9490C (.Z(FE_OFN70_g9490C),.A(g9490C));
BUF_X3 FE_OFC69_g9392C (.Z(FE_OFN69_g9392C),.A(FE_OFN68_g9392C));
BUF_X3 FE_OFC68_g9392C (.Z(FE_OFN68_g9392C),.A(g9392C));
BUF_X3 FE_OFC67_g9367C (.Z(FE_OFN67_g9367C),.A(g9367C));
BUF_X3 FE_OFC64_g9536C (.Z(FE_OFN64_g9536C),.A(g9536C));
BUF_X3 FE_OFC63_g9474C (.Z(FE_OFN63_g9474C),.A(g9474C));
BUF_X3 FE_OFC62_g9274C (.Z(FE_OFN62_g9274C),.A(g9274C));
BUF_X3 FE_OFC61_g9624C (.Z(FE_OFN61_g9624C),.A(FE_OFN60_g9624C));
BUF_X3 FE_OFC60_g9624C (.Z(FE_OFN60_g9624C),.A(g9624C));
INV_X1 FE_OFC59_g9432C (.ZN(FE_OFN59_g9432C),.A(FE_OFN57_g9432C));
INV_X1 FE_OFC57_g9432C (.ZN(FE_OFN57_g9432C),.A(g9432C));
BUF_X3 FE_OFC56_g9052C (.Z(FE_OFN56_g9052C),.A(FE_OFN54_g9052C));
BUF_X3 FE_OFC54_g9052C (.Z(FE_OFN54_g9052C),.A(g9052C));
BUF_X3 FE_OFC53_g9173C (.Z(FE_OFN53_g9173C),.A(FE_OFN52_g9173C));
BUF_X3 FE_OFC52_g9173C (.Z(FE_OFN52_g9173C),.A(g9173C));
BUF_X3 FE_OFC51_g9111C (.Z(FE_OFN51_g9111C),.A(g9111C));
BUF_X3 FE_OFC50_g9030C (.Z(FE_OFN50_g9030C),.A(FE_OFN49_g9030C));
BUF_X3 FE_OFC49_g9030C (.Z(FE_OFN49_g9030C),.A(g9030C));
BUF_X3 FE_OFC48_g9151C (.Z(FE_OFN48_g9151C),.A(FE_OFN47_g9151C));
BUF_X3 FE_OFC47_g9151C (.Z(FE_OFN47_g9151C),.A(g9151C));
BUF_X3 FE_OFC46_g9125C (.Z(FE_OFN46_g9125C),.A(FE_OFN45_g9125C));
BUF_X3 FE_OFC45_g9125C (.Z(FE_OFN45_g9125C),.A(FE_OFN44_g9125C));
BUF_X3 FE_OFC44_g9125C (.Z(FE_OFN44_g9125C),.A(g9125C));
BUF_X3 FE_OFC42_g9205C (.Z(FE_OFN42_g9205C),.A(g9205C));
BUF_X3 FE_OFC40_g9240C (.Z(FE_OFN40_g9240C),.A(g9240C));
BUF_X3 FE_OFC39_g9223C (.Z(FE_OFN39_g9223C),.A(g9223C));
BUF_X3 FE_OFC35_g9785C (.Z(FE_OFN35_g9785C),.A(FE_OFN34_g9785C));
BUF_X3 FE_OFC34_g9785C (.Z(FE_OFN34_g9785C),.A(g9785C));
BUF_X3 FE_OFC33_g9454C (.Z(FE_OFN33_g9454C),.A(FE_OFN32_g9454C));
BUF_X3 FE_OFC32_g9454C (.Z(FE_OFN32_g9454C),.A(g9454C));
BUF_X3 FE_OFC27_g11519C (.Z(FE_OFN27_g11519C),.A(g11519C));
BUF_X3 FE_OFC21_g10702C (.Z(FE_OFN21_g10702C),.A(FE_OFN20_g10702C));
BUF_X3 FE_OFC20_g10702C (.Z(FE_OFN20_g10702C),.A(FE_OFN18_g10702C));
BUF_X3 FE_OFC18_g10702C (.Z(FE_OFN18_g10702C),.A(FE_OFN13_g10702C));
INV_X1 FE_OFC17_g10702C (.ZN(FE_OFN17_g10702C),.A(FE_OFN15_g10702C));
INV_X1 FE_OFC15_g10702C (.ZN(FE_OFN15_g10702C),.A(FE_OFN14_g10702C));
BUF_X3 FE_OFC14_g10702C (.Z(FE_OFN14_g10702C),.A(FE_OFN9_g10702C));
INV_X1 FE_OFC13_g10702C (.ZN(FE_OFN13_g10702C),.A(FE_OFN10_g10702C));
INV_X1 FE_OFC10_g10702C (.ZN(FE_OFN10_g10702C),.A(FE_OFN9_g10702C));
BUF_X3 FE_OFC9_g10702C (.Z(FE_OFN9_g10702C),.A(FE_OFN8_g10702C));
BUF_X3 FE_OFC8_g10702C (.Z(FE_OFN8_g10702C),.A(FE_OFN7_g10702C));
BUF_X3 FE_OFC7_g10702C (.Z(FE_OFN7_g10702C),.A(g10702C));
BUF_X3 FE_OFC4_g10950C (.Z(FE_OFN4_g10950C),.A(FE_OFN3_g10950C));
INV_X1 FE_OFC3_g10950C (.ZN(FE_OFN3_g10950C),.A(FE_OFN0_g10950C));
INV_X1 FE_OFC0_g10950C (.ZN(FE_OFN0_g10950C),.A(g10950C));
INV_X1 U_g2299C (.ZN(g2299C),.A(g1707C));
INV_X1 U_g9291C (.ZN(g9291C),.A(FE_OFN79_g8700C));
INV_X4 U_I7048C (.ZN(I7048C),.A(g2807C));
INV_X1 U_g1981C (.ZN(g1981C),.A(g650C));
INV_X1 U_g3982C (.ZN(g3982C),.A(g2118C));
INV_X1 U_g3629C (.ZN(g3629C),.A(FE_OFN266_g18C));
INV_X1 U_g6842C (.ZN(g6842C),.A(I9769C));
INV_X1 U_g8617C (.ZN(g8617C),.A(g8465C));
INV_X1 U_g2078C (.ZN(g2078C),.A(g135C));
INV_X1 U_g2340C (.ZN(g2340C),.A(g1918C));
INV_X1 U_g7684C (.ZN(g7684C),.A(FE_OFN83_g2176C));
INV_X1 U_g3800C (.ZN(g3800C),.A(FE_OFN250_g471C));
INV_X1 U_g6941C (.ZN(g6941C),.A(FE_OFN88_g2178C));
INV_X1 U_g2435C (.ZN(g2435C),.A(g201C));
INV_X4 U_g4010C (.ZN(g4010C),.A(g3744C));
INV_X1 U_g2082C (.ZN(g2082C),.A(g1371C));
INV_X1 U_g5519C (.ZN(g5519C),.A(g4811C));
INV_X1 U_g10668C (.ZN(g10668C),.A(g10563C));
INV_X1 U_g4172C (.ZN(g4172C),.A(g2057C));
INV_X1 U_g8709C (.ZN(g8709C),.A(g8451C));
INV_X1 U_g2214C (.ZN(g2214C),.A(g115C));
INV_X1 U_I7847C (.ZN(I7847C),.A(g3435C));
INV_X1 U_g8340C (.ZN(g8340C),.A(I13400C));
INV_X1 U_g4566C (.ZN(g4566C),.A(g3753C));
INV_X1 U_g3348C (.ZN(g3348C),.A(FE_OFN267_g109C));
INV_X1 U_I15968C (.ZN(I15968C),.A(g10408C));
INV_X1 U_g11060C (.ZN(g11060C),.A(g10937C));
INV_X1 U_I15855C (.ZN(I15855C),.A(g10336C));
INV_X1 U_g6270C (.ZN(g6270C),.A(I9383C));
INV_X1 U_g10679C (.ZN(g10679C),.A(g10584C));
INV_X1 U_g1968C (.ZN(g1968C),.A(g369C));
INV_X1 U_g5659C (.ZN(g5659C),.A(I7771C));
INV_X1 U_I15503C (.ZN(I15503C),.A(g9995C));
INV_X1 U_g8110C (.ZN(g8110C),.A(g7996C));
INV_X1 U_g2556C (.ZN(g2556C),.A(g186C));
INV_X1 U_I7817C (.ZN(I7817C),.A(g3399C));
INV_X1 U_g2222C (.ZN(g2222C),.A(g158C));
INV_X1 U_I13373C (.ZN(I13373C),.A(g8226C));
INV_X1 U_g4202C (.ZN(g4202C),.A(I5430C));
INV_X1 U_I9880C (.ZN(I9880C),.A(g5405C));
INV_X1 U_g4094C (.ZN(g4094C),.A(g2744C));
INV_X1 U_g4567C (.ZN(g4567C),.A(g3374C));
INV_X1 U_I14312C (.ZN(I14312C),.A(g8814C));
INV_X1 U_g11111C (.ZN(g11111C),.A(g10702C));
INV_X1 U_g4776C (.ZN(g4776C),.A(FE_OFN344_g3586C));
INV_X1 U_I15986C (.ZN(I15986C),.A(g10417C));
INV_X1 U_g2237C (.ZN(g2237C),.A(g713C));
INV_X1 U_g7897C (.ZN(g7897C),.A(g7712C));
INV_X1 U_g3121C (.ZN(g3121C),.A(FE_OFN352_g109C));
INV_X1 U_g5420C (.ZN(g5420C),.A(g4300C));
INV_X1 U_g10455C (.ZN(g10455C),.A(I15956C));
INV_X1 U_g2557C (.ZN(g2557C),.A(g1840C));
INV_X1 U_g9097C (.ZN(g9097C),.A(g8700C));
INV_X1 U_g3938C (.ZN(g3938C),.A(g2299C));
INV_X1 U_g8563C (.ZN(g8563C),.A(I7829C));
INV_X1 U_g6259C (.ZN(g6259C),.A(g2175C));
INV_X1 U_g4179C (.ZN(g4179C),.A(g1992C));
INV_X1 U_g7682C (.ZN(g7682C),.A(FE_OFN83_g2176C));
INV_X1 U_g4379C (.ZN(g4379C),.A(g3698C));
INV_X1 U_I4917C (.ZN(I4917C),.A(g584C));
INV_X1 U_g2254C (.ZN(g2254C),.A(g131C));
INV_X1 U_g4289C (.ZN(g4289C),.A(FE_OFN298_g3015C));
INV_X1 U_g4777C (.ZN(g4777C),.A(g3992C));
INV_X1 U_g8089C (.ZN(g8089C),.A(g7934C));
INV_X1 U_g2438C (.ZN(g2438C),.A(g243C));
INV_X1 U_g4271C (.ZN(g4271C),.A(g2024C));
INV_X1 U_g7045C (.ZN(g7045C),.A(g6003C));
INV_X1 U_I5424C (.ZN(I5424C),.A(g910C));
INV_X1 U_g2212C (.ZN(g2212C),.A(g686C));
INV_X1 U_g3141C (.ZN(g3141C),.A(g2563C));
INV_X1 U_g3710C (.ZN(g3710C),.A(g3215C));
INV_X1 U_g7920C (.ZN(g7920C),.A(g7516C));
INV_X1 U_g2229C (.ZN(g2229C),.A(g162C));
INV_X1 U_I15157C (.ZN(I15157C),.A(g9931C));
INV_X1 U_g11157C (.ZN(g11157C),.A(FE_OFN3_g10950C));
INV_X1 U_g4209C (.ZN(g4209C),.A(I5002C));
INV_X1 U_I9279C (.ZN(I9279C),.A(g91C));
INV_X1 U_I5044C (.ZN(I5044C),.A(g1182C));
INV_X1 U_I15287C (.ZN(I15287C),.A(g9968C));
INV_X1 U_g2249C (.ZN(g2249C),.A(g127C));
INV_X1 U_g11596C (.ZN(g11596C),.A(g11580C));
INV_X1 U_g11243C (.ZN(g11243C),.A(FE_OFN8_g10702C));
INV_X1 U_g6266C (.ZN(g6266C),.A(g2208C));
INV_X1 U_g8062C (.ZN(g8062C),.A(I4783C));
INV_X1 U_I5414C (.ZN(I5414C),.A(g904C));
INV_X1 U_g3628C (.ZN(g3628C),.A(g3111C));
INV_X1 U_g6255C (.ZN(g6255C),.A(I9237C));
INV_X1 U_g4175C (.ZN(g4175C),.A(g1988C));
INV_X1 U_g6081C (.ZN(g6081C),.A(g4977C));
INV_X1 U_g7910C (.ZN(g7910C),.A(g7460C));
INV_X1 U_g4285C (.ZN(g4285C),.A(g3688C));
INV_X1 U_g6354C (.ZN(g6354C),.A(g5867C));
INV_X1 U_g2031C (.ZN(g2031C),.A(g1690C));
INV_X1 U_g8085C (.ZN(g8085C),.A(g7932C));
INV_X1 U_g2176C (.ZN(g2176C),.A(g82C));
INV_X1 U_g7883C (.ZN(g7883C),.A(g7246C));
INV_X1 U_g4737C (.ZN(g4737C),.A(g3440C));
INV_X1 U_I13351C (.ZN(I13351C),.A(g8214C));
INV_X1 U_g6267C (.ZN(g6267C),.A(I9326C));
INV_X1 U_g3440C (.ZN(g3440C),.A(g3041C));
INV_X1 U_g2610C (.ZN(g2610C),.A(I4917C));
INV_X1 U_g4205C (.ZN(g4205C),.A(I4992C));
INV_X1 U_g10883C (.ZN(g10883C),.A(g10809C));
INV_X1 U_g5521C (.ZN(g5521C),.A(FE_OFN221_g3440C));
INV_X1 U_I6260C (.ZN(I6260C),.A(g1696C));
INV_X1 U_I9311C (.ZN(I9311C),.A(g103C));
INV_X1 U_I5579C (.ZN(I5579C),.A(g1197C));
INV_X1 U_g10439C (.ZN(g10439C),.A(g10334C));
INV_X1 U_g5878C (.ZN(g5878C),.A(g5309C));
INV_X1 U_g6932C (.ZN(g6932C),.A(I7829C));
INV_X1 U_g4273C (.ZN(g4273C),.A(FE_OFN133_g3015C));
INV_X1 U_g5658C (.ZN(g5658C),.A(I7752C));
INV_X1 U_g7467C (.ZN(g7467C),.A(FE_OFN84_g2176C));
INV_X1 U_g1990C (.ZN(g1990C),.A(g774C));
INV_X1 U_I13436C (.ZN(I13436C),.A(g8187C));
INV_X1 U_g2399C (.ZN(g2399C),.A(g605C));
INV_X1 U_g8980C (.ZN(g8980C),.A(I14306C));
INV_X1 U_g6716C (.ZN(g6716C),.A(FE_OFN115_g4807C));
INV_X1 U_g7685C (.ZN(g7685C),.A(FE_OFN87_g2176C));
INV_X1 U_g8849C (.ZN(g8849C),.A(g8745C));
INV_X1 U_I7840C (.ZN(I7840C),.A(g3431C));
INV_X1 U_g10852C (.ZN(g10852C),.A(g10739C));
INV_X1 U_g7562C (.ZN(g7562C),.A(FE_OFN91_g2172C));
INV_X1 U_g6258C (.ZN(g6258C),.A(g2172C));
INV_X1 U_g4178C (.ZN(g4178C),.A(g1991C));
INV_X4 U_g4679C (.ZN(g4679C),.A(FE_OFN293_g3015C));
INV_X1 U_g3776C (.ZN(g3776C),.A(g2579C));
INV_X1 U_g2008C (.ZN(g2008C),.A(g971C));
INV_X1 U_g6274C (.ZN(g6274C),.A(I9293C));
INV_X1 U_g2336C (.ZN(g2336C),.A(g1900C));
INV_X1 U_g3521C (.ZN(g3521C),.A(FE_OFN359_g18C));
INV_X1 U_g6280C (.ZN(g6280C),.A(g2253C));
INV_X1 U_I6962C (.ZN(I6962C),.A(g2791C));
INV_X1 U_g2230C (.ZN(g2230C),.A(g704C));
INV_X1 U_g4437C (.ZN(g4437C),.A(FE_OFN235_g2024C));
INV_X1 U_g4208C (.ZN(g4208C),.A(I5588C));
INV_X1 U_g7505C (.ZN(g7505C),.A(FE_OFN87_g2176C));
INV_X1 U_I15974C (.ZN(I15974C),.A(g10411C));
INV_X1 U_g2550C (.ZN(g2550C),.A(g1834C));
INV_X1 U_g10400C (.ZN(g10400C),.A(g10348C));
INV_X1 U_I9282C (.ZN(I9282C),.A(g101C));
INV_X1 U_I5584C (.ZN(I5584C),.A(g1200C));
INV_X4 U_g9490C (.ZN(g9490C),.A(g9324C));
INV_X1 U_g2395C (.ZN(g2395C),.A(g231C));
INV_X1 U_g8465C (.ZN(g8465C),.A(g8289C));
INV_X1 U_g6403C (.ZN(g6403C),.A(g5013C));
INV_X1 U_I15510C (.ZN(I15510C),.A(g10013C));
INV_X1 U_g2248C (.ZN(g2248C),.A(g99C));
INV_X1 U_g3744C (.ZN(g3744C),.A(FE_OFN269_g109C));
INV_X1 U_I4883C (.ZN(I4883C),.A(g581C));
INV_X1 U_g7688C (.ZN(g7688C),.A(FE_OFN83_g2176C));
INV_X1 U_g2481C (.ZN(g2481C),.A(g882C));
INV_X1 U_g10683C (.ZN(g10683C),.A(g10385C));
INV_X1 U_I5070C (.ZN(I5070C),.A(g1194C));
INV_X1 U_g4888C (.ZN(g4888C),.A(I5101C));
INV_X1 U_g4171C (.ZN(g4171C),.A(I6962C));
INV_X1 U_g4787C (.ZN(g4787C),.A(g3423C));
INV_X1 U_g6447C (.ZN(g6447C),.A(FE_OFN218_g5557C));
INV_X1 U_g3092C (.ZN(g3092C),.A(g639C));
INV_X1 U_g4281C (.ZN(g4281C),.A(g3586C));
INV_X1 U_g5613C (.ZN(g5613C),.A(FE_OFN131_g3015C));
INV_X1 U_g8255C (.ZN(g8255C),.A(g7986C));
INV_X1 U_g8081C (.ZN(g8081C),.A(g8000C));
INV_X1 U_I5406C (.ZN(I5406C),.A(g898C));
INV_X1 U_I4780C (.ZN(I4780C),.A(g872C));
INV_X1 U_g10584C (.ZN(g10584C),.A(g10522C));
INV_X1 U_g6272C (.ZN(g6272C),.A(I9268C));
INV_X1 U_g8783C (.ZN(g8783C),.A(g8746C));
INV_X1 U_g8979C (.ZN(g8979C),.A(I14303C));
INV_X1 U_g4201C (.ZN(g4201C),.A(I5427C));
INV_X1 U_I5445C (.ZN(I5445C),.A(g922C));
INV_X1 U_g4449C (.ZN(g4449C),.A(g4144C));
INV_X1 U_g7696C (.ZN(g7696C),.A(FE_OFN86_g2176C));
INV_X1 U_g8828C (.ZN(g8828C),.A(g8744C));
INV_X1 U_g2677C (.ZN(g2677C),.A(g2034C));
INV_X1 U_g10361C (.ZN(g10361C),.A(g10268C));
INV_X1 U_g3737C (.ZN(g3737C),.A(g2506C));
INV_X1 U_I9332C (.ZN(I9332C),.A(g104C));
INV_X1 U_g9525C (.ZN(g9525C),.A(g9257C));
INV_X1 U_g2198C (.ZN(g2198C),.A(g668C));
INV_X1 U_I7771C (.ZN(I7771C),.A(g3418C));
INV_X1 U_g3523C (.ZN(g3523C),.A(g1845C));
INV_X1 U_g2241C (.ZN(g2241C),.A(g722C));
INV_X1 U_g7681C (.ZN(g7681C),.A(FE_OFN87_g2176C));
INV_X1 U_g7697C (.ZN(g7697C),.A(g7101C));
INV_X1 U_g7914C (.ZN(g7914C),.A(g7651C));
INV_X1 U_g8349C (.ZN(g8349C),.A(I13427C));
INV_X1 U_g6260C (.ZN(g6260C),.A(g2178C));
INV_X1 U_I14319C (.ZN(I14319C),.A(g8816C));
INV_X1 U_g10463C (.ZN(g10463C),.A(I15980C));
INV_X1 U_I5388C (.ZN(I5388C),.A(g889C));
INV_X1 U_g2211C (.ZN(g2211C),.A(g153C));
INV_X1 U_g6279C (.ZN(g6279C),.A(g2248C));
INV_X1 U_g3983C (.ZN(g3983C),.A(g3222C));
INV_X1 U_I5430C (.ZN(I5430C),.A(g916C));
INV_X4 U_g4678C (.ZN(g4678C),.A(g3546C));
INV_X1 U_g3543C (.ZN(g3543C),.A(g3101C));
INV_X1 U_g9507C (.ZN(g9507C),.A(g9268C));
INV_X1 U_g10421C (.ZN(g10421C),.A(g10331C));
INV_X1 U_g8352C (.ZN(g8352C),.A(I13436C));
INV_X1 U_g7460C (.ZN(g7460C),.A(FE_OFN85_g2176C));
INV_X1 U_g2083C (.ZN(g2083C),.A(g139C));
INV_X1 U_I6360C (.ZN(I6360C),.A(g1713C));
INV_X1 U_I4992C (.ZN(I4992C),.A(g1170C));
INV_X1 U_I16982C (.ZN(I16982C),.A(g10629C));
INV_X1 U_g8599C (.ZN(g8599C),.A(g8546C));
INV_X1 U_g6253C (.ZN(g6253C),.A(I9479C));
INV_X1 U_g2061C (.ZN(g2061C),.A(g1828C));
INV_X1 U_g2187C (.ZN(g2187C),.A(g746C));
INV_X1 U_g4173C (.ZN(g4173C),.A(g1984C));
INV_X1 U_g8984C (.ZN(g8984C),.A(I14319C));
INV_X1 U_g2446C (.ZN(g2446C),.A(g1400C));
INV_X1 U_g11575C (.ZN(g11575C),.A(g11561C));
INV_X1 U_g2345C (.ZN(g2345C),.A(g1936C));
INV_X1 U_g8106C (.ZN(g8106C),.A(g7950C));
INV_X1 U_g6586C (.ZN(g6586C),.A(FE_OFN118_g4807C));
INV_X1 U_g8061C (.ZN(g8061C),.A(I4780C));
INV_X1 U_g5808C (.ZN(g5808C),.A(g85C));
INV_X1 U_I5418C (.ZN(I5418C),.A(g907C));
INV_X1 U_g4203C (.ZN(g4203C),.A(I5441C));
INV_X1 U_g2016C (.ZN(g2016C),.A(g1361C));
INV_X1 U_I16252C (.ZN(I16252C),.A(g10515C));
INV_X1 U_I9273C (.ZN(I9273C),.A(g47C));
INV_X1 U_g2251C (.ZN(g2251C),.A(g731C));
INV_X1 U_g2047C (.ZN(g2047C),.A(g1857C));
INV_X1 U_g10927C (.ZN(g10927C),.A(FE_OFN17_g10702C));
INV_X1 U_g6275C (.ZN(g6275C),.A(I9308C));
INV_X1 U_g4216C (.ZN(g4216C),.A(I5070C));
INV_X1 U_g8858C (.ZN(g8858C),.A(g8743C));
INV_X1 U_g4671C (.ZN(g4671C),.A(g3354C));
INV_X1 U_g8115C (.ZN(g8115C),.A(g7953C));
INV_X1 U_g2612C (.ZN(g2612C),.A(I4948C));
INV_X1 U_g2017C (.ZN(g2017C),.A(g1218C));
INV_X1 U_g6284C (.ZN(g6284C),.A(I9332C));
INV_X1 U_g7683C (.ZN(g7683C),.A(FE_OFN87_g2176C));
INV_X1 U_I5101C (.ZN(I5101C),.A(g1960C));
INV_X1 U_g2328C (.ZN(g2328C),.A(g1882C));
INV_X1 U_g2542C (.ZN(g2542C),.A(g1868C));
INV_X1 U_g2330C (.ZN(g2330C),.A(g1891C));
INV_X1 U_g7949C (.ZN(g7949C),.A(FE_OFN211_g7246C));
INV_X1 U_I5041C (.ZN(I5041C),.A(g1179C));
INV_X1 U_g1992C (.ZN(g1992C),.A(g782C));
INV_X1 U_g8978C (.ZN(g8978C),.A(I14299C));
INV_X1 U_I5441C (.ZN(I5441C),.A(g919C));
INV_X1 U_g4365C (.ZN(g4365C),.A(g3880C));
INV_X1 U_g8982C (.ZN(g8982C),.A(I14312C));
INV_X1 U_g8234C (.ZN(g8234C),.A(FE_OFN198_g7697C));
INV_X1 U_g8328C (.ZN(g8328C),.A(I13364C));
INV_X1 U_g4196C (.ZN(g4196C),.A(I5245C));
INV_X1 U_g2456C (.ZN(g2456C),.A(g1397C));
INV_X1 U_g7919C (.ZN(g7919C),.A(g7512C));
INV_X1 U_g5105C (.ZN(g5105C),.A(I4783C));
INV_X1 U_g1976C (.ZN(g1976C),.A(g643C));
INV_X1 U_g7952C (.ZN(g7952C),.A(FE_OFN210_g7246C));
INV_X1 U_I4820C (.ZN(I4820C),.A(g865C));
INV_X1 U_g2355C (.ZN(g2355C),.A(I5435C));
INV_X1 U_I14315C (.ZN(I14315C),.A(g8815C));
INV_X1 U_g4467C (.ZN(g4467C),.A(g3829C));
INV_X1 U_g4290C (.ZN(g4290C),.A(FE_OFN102_g3586C));
INV_X1 U_g7527C (.ZN(g7527C),.A(FE_OFN85_g2176C));
INV_X1 U_I9265C (.ZN(I9265C),.A(g46C));
INV_X1 U_g8056C (.ZN(g8056C),.A(g7671C));
INV_X1 U_g4181C (.ZN(g4181C),.A(g2449C));
INV_X1 U_g4381C (.ZN(g4381C),.A(FE_OFN296_g3914C));
INV_X1 U_g2118C (.ZN(g2118C),.A(g1854C));
INV_X1 U_I6273C (.ZN(I6273C),.A(FE_OFN363_I5565C));
INV_X1 U_g10629C (.ZN(g10629C),.A(g10583C));
INV_X1 U_g4197C (.ZN(g4197C),.A(I5410C));
INV_X1 U_g2652C (.ZN(g2652C),.A(g2008C));
INV_X1 U_g2057C (.ZN(g2057C),.A(g754C));
INV_X1 U_g10628C (.ZN(g10628C),.A(I16252C));
INV_X1 U_g3539C (.ZN(g3539C),.A(g3015C));
INV_X1 U_g4263C (.ZN(g4263C),.A(FE_OFN103_g3586C));
INV_X1 U_I9296C (.ZN(I9296C),.A(g102C));
INV_X1 U_I13323C (.ZN(I13323C),.A(g8203C));
INV_X1 U_g2549C (.ZN(g2549C),.A(g1386C));
INV_X1 U_g6278C (.ZN(g6278C),.A(I9371C));
INV_X1 U_g5261C (.ZN(g5261C),.A(g4640C));
INV_X1 U_g3419C (.ZN(g3419C),.A(g3104C));
INV_X1 U_I7829C (.ZN(I7829C),.A(g3425C));
INV_X1 U_g7516C (.ZN(g7516C),.A(FE_OFN82_g2176C));
INV_X1 U_g6282C (.ZN(g6282C),.A(I9296C));
INV_X1 U_g9802C (.ZN(g9802C),.A(g9490C));
INV_X1 U_g8318C (.ZN(g8318C),.A(I13338C));
INV_X1 U_g3086C (.ZN(g3086C),.A(g2276C));
INV_X1 U_g2253C (.ZN(g2253C),.A(g100C));
INV_X1 U_I9371C (.ZN(I9371C),.A(g96C));
INV_X1 U_I5383C (.ZN(I5383C),.A(g886C));
INV_X1 U_g2606C (.ZN(g2606C),.A(I4876C));
INV_X1 U_I5588C (.ZN(I5588C),.A(g1203C));
INV_X1 U_g7907C (.ZN(g7907C),.A(g7664C));
INV_X1 U_g4673C (.ZN(g4673C),.A(FE_OFN348_g3015C));
INV_X1 U_g2570C (.ZN(g2570C),.A(g207C));
INV_X1 U_g7915C (.ZN(g7915C),.A(g7473C));
INV_X1 U_g10377C (.ZN(g10377C),.A(I15855C));
INV_X1 U_g6264C (.ZN(g6264C),.A(g2176C));
INV_X1 U_g2607C (.ZN(g2607C),.A(I4883C));
INV_X1 U_g2506C (.ZN(g2506C),.A(g636C));
INV_X1 U_I16717C (.ZN(I16717C),.A(g10779C));
INV_X1 U_g3491C (.ZN(g3491C),.A(g1107C));
INV_X1 U_I7852C (.ZN(I7852C),.A(g3438C));
INV_X1 U_g2275C (.ZN(g2275C),.A(g757C));
INV_X1 U_g3007C (.ZN(g3007C),.A(I6240C));
INV_X1 U_g2374C (.ZN(g2374C),.A(g591C));
INV_X1 U_I9268C (.ZN(I9268C),.A(g90C));
INV_X1 U_g9424C (.ZN(g9424C),.A(g9291C));
INV_X1 U_g6271C (.ZN(g6271C),.A(I9259C));
INV_X1 U_g3793C (.ZN(g3793C),.A(FE_OFN248_g466C));
INV_X1 U_I7825C (.ZN(I7825C),.A(g3414C));
INV_X1 U_g2420C (.ZN(g2420C),.A(g237C));
INV_X1 U_g3664C (.ZN(g3664C),.A(g3209C));
INV_X1 U_g5509C (.ZN(g5509C),.A(g4739C));
INV_X1 U_g8985C (.ZN(g8985C),.A(I14326C));
INV_X1 U_g4608C (.ZN(g4608C),.A(FE_OFN141_g3829C));
INV_X1 U_g5816C (.ZN(g5816C),.A(g1810C));
INV_X1 U_I5060C (.ZN(I5060C),.A(g1191C));
INV_X1 U_I14306C (.ZN(I14306C),.A(g8812C));
INV_X1 U_g9961C (.ZN(g9961C),.A(I15157C));
INV_X1 U_g7438C (.ZN(g7438C),.A(FE_OFN195_g6488C));
INV_X1 U_g8100C (.ZN(g8100C),.A(g7947C));
INV_X1 U_g5101C (.ZN(g5101C),.A(I4780C));
INV_X1 U_g7918C (.ZN(g7918C),.A(g7505C));
INV_X1 U_g6262C (.ZN(g6262C),.A(I9273C));
INV_X1 U_g2648C (.ZN(g2648C),.A(I4820C));
INV_X1 U_g2410C (.ZN(g2410C),.A(g1453C));
INV_X1 U_g8323C (.ZN(g8323C),.A(I13351C));
INV_X1 U_I5053C (.ZN(I5053C),.A(g1188C));
INV_X1 U_g6285C (.ZN(g6285C),.A(I9352C));
INV_X1 U_g2172C (.ZN(g2172C),.A(g43C));
INV_X1 U_I13364C (.ZN(I13364C),.A(g8221C));
INV_X1 U_g2343C (.ZN(g2343C),.A(g1927C));
INV_X1 U_g4210C (.ZN(g4210C),.A(I5020C));
INV_X1 U_I4876C (.ZN(I4876C),.A(g580C));
INV_X1 U_g8566C (.ZN(g8566C),.A(I7852C));
INV_X1 U_g2202C (.ZN(g2202C),.A(g148C));
INV_X1 U_g6926C (.ZN(g6926C),.A(I7825C));
INV_X1 U_g8548C (.ZN(g8548C),.A(g8390C));
INV_X1 U_g2518C (.ZN(g2518C),.A(g590C));
INV_X1 U_g6273C (.ZN(g6273C),.A(I9279C));
INV_X1 U_g10801C (.ZN(g10801C),.A(I16507C));
INV_X1 U_g4739C (.ZN(g4739C),.A(g4117C));
INV_X1 U_g6269C (.ZN(g6269C),.A(I9368C));
INV_X1 U_g8313C (.ZN(g8313C),.A(I13323C));
INV_X1 U_I9308C (.ZN(I9308C),.A(g93C));
INV_X1 U_g4294C (.ZN(g4294C),.A(g3664C));
INV_X1 U_g3723C (.ZN(g3723C),.A(g3071C));
INV_X1 U_g10457C (.ZN(g10457C),.A(I15962C));
INV_X1 U_g8094C (.ZN(g8094C),.A(g7987C));
INV_X1 U_g2050C (.ZN(g2050C),.A(g1861C));
INV_X1 U_g7473C (.ZN(g7473C),.A(FE_OFN87_g2176C));
INV_X1 U_g2777C (.ZN(g2777C),.A(FE_OFN224_g2276C));
INV_X1 U_g2271C (.ZN(g2271C),.A(g877C));
INV_X1 U_g2611C (.ZN(g2611C),.A(I4935C));
INV_X1 U_g3368C (.ZN(g3368C),.A(g2459C));
INV_X1 U_g1987C (.ZN(g1987C),.A(g762C));
INV_X4 U_I8869C (.ZN(I8869C),.A(g4421C));
INV_X1 U_I9290C (.ZN(I9290C),.A(FE_OFN277_g48C));
INV_X1 U_I4948C (.ZN(I4948C),.A(g586C));
INV_X1 U_g8271C (.ZN(g8271C),.A(g1810C));
INV_X1 U_g1991C (.ZN(g1991C),.A(g778C));
INV_X1 U_g11199C (.ZN(g11199C),.A(FE_OFN21_g10702C));
INV_X1 U_g8981C (.ZN(g8981C),.A(I14309C));
INV_X1 U_I15365C (.ZN(I15365C),.A(g10025C));
INV_X1 U_g7852C (.ZN(g7852C),.A(FE_OFN209_g6863C));
INV_X1 U_g7923C (.ZN(g7923C),.A(g7527C));
INV_X1 U_g10431C (.ZN(g10431C),.A(g10328C));
INV_X1 U_g6265C (.ZN(g6265C),.A(I9276C));
INV_X1 U_g4782C (.ZN(g4782C),.A(g4089C));
INV_X1 U_g4292C (.ZN(g4292C),.A(FE_OFN136_g3863C));
INV_X1 U_g3760C (.ZN(g3760C),.A(g3003C));
INV_X1 U_I5435C (.ZN(I5435C),.A(g18C));
INV_X1 U_g5117C (.ZN(g5117C),.A(FE_OFN144_g4682C));
INV_X4 U_g2175C (.ZN(g2175C),.A(g44C));
INV_X1 U_I9368C (.ZN(I9368C),.A(g87C));
INV_X4 U_g2024C (.ZN(g2024C),.A(g1718C));
INV_X1 U_g6281C (.ZN(g6281C),.A(I9282C));
INV_X1 U_g3327C (.ZN(g3327C),.A(g23C));
INV_X4 U_g2424C (.ZN(g2424C),.A(FE_OFN241_g1690C));
INV_X1 U_I5002C (.ZN(I5002C),.A(g1173C));
INV_X1 U_g7550C (.ZN(g7550C),.A(FE_OFN96_g2169C));
INV_X1 U_g2077C (.ZN(g2077C),.A(g219C));
INV_X1 U_g3103C (.ZN(g3103C),.A(g1212C));
INV_X1 U_g7913C (.ZN(g7913C),.A(g7467C));
INV_X1 U_g6109C (.ZN(g6109C),.A(g48C));
INV_X1 U_g6449C (.ZN(g6449C),.A(g5557C));
INV_X1 U_g2273C (.ZN(g2273C),.A(g881C));
INV_X1 U_g7692C (.ZN(g7692C),.A(g2176C));
INV_X1 U_g7497C (.ZN(g7497C),.A(FE_OFN85_g2176C));
INV_X1 U_g2444C (.ZN(g2444C),.A(g876C));
INV_X1 U_g8099C (.ZN(g8099C),.A(g7990C));
INV_X1 U_I9326C (.ZN(I9326C),.A(FE_OFN271_g85C));
INV_X1 U_g6268C (.ZN(g6268C),.A(I9346C));
INV_X1 U_g10676C (.ZN(g10676C),.A(g10570C));
INV_X1 U_g1993C (.ZN(g1993C),.A(g786C));
INV_X1 U_I9383C (.ZN(I9383C),.A(g88C));
INV_X1 U_g8983C (.ZN(g8983C),.A(I14315C));
INV_X1 U_I5254C (.ZN(I5254C),.A(g1700C));
INV_X1 U_I14303C (.ZN(I14303C),.A(g8811C));
INV_X1 U_g2178C (.ZN(g2178C),.A(g45C));
INV_X1 U_I4900C (.ZN(I4900C),.A(g583C));
INV_X1 U_g3060C (.ZN(g3060C),.A(FE_OFN245_g1690C));
INV_X1 U_g4214C (.ZN(g4214C),.A(I5053C));
INV_X1 U_I9346C (.ZN(I9346C),.A(g86C));
INV_X1 U_g2382C (.ZN(g2382C),.A(g599C));
INV_X1 U_g3784C (.ZN(g3784C),.A(FE_OFN254_g461C));
INV_X1 U_I17413C (.ZN(I17413C),.A(g11425C));
INV_X1 U_g7677C (.ZN(g7677C),.A(FE_OFN85_g2176C));
INV_X4 U_g4002C (.ZN(g4002C),.A(FE_OFN155_g3121C));
INV_X1 U_g3479C (.ZN(g3479C),.A(g1101C));
INV_X1 U_g11489C (.ZN(g11489C),.A(I17413C));
INV_X1 U_g6131C (.ZN(g6131C),.A(g5548C));
INV_X1 U_g3390C (.ZN(g3390C),.A(g2045C));
INV_X1 U_g5627C (.ZN(g5627C),.A(FE_OFN132_g3015C));
INV_X1 U_g3501C (.ZN(g3501C),.A(FE_OFN240_g1110C));
INV_X1 U_g8335C (.ZN(g8335C),.A(I13385C));
INV_X1 U_g2095C (.ZN(g2095C),.A(g143C));
INV_X1 U_g2208C (.ZN(g2208C),.A(g84C));
INV_X1 U_g2579C (.ZN(g2579C),.A(g1969C));
INV_X1 U_I14326C (.ZN(I14326C),.A(g8818C));
INV_X1 U_g6283C (.ZN(g6283C),.A(I9311C));
INV_X1 U_g6920C (.ZN(g6920C),.A(I7817C));
INV_X1 U_g8095C (.ZN(g8095C),.A(g7942C));
INV_X1 U_g6718C (.ZN(g6718C),.A(FE_OFN116_g4807C));
INV_X1 U_g2364C (.ZN(g2364C),.A(g611C));
INV_X1 U_g4194C (.ZN(g4194C),.A(I5399C));
INV_X1 U_g2054C (.ZN(g2054C),.A(g1864C));
INV_X1 U_g6261C (.ZN(g6261C),.A(I9265C));
INV_X1 U_g2725C (.ZN(g2725C),.A(g2018C));
INV_X1 U_g5503C (.ZN(g5503C),.A(FE_OFN204_g3664C));
INV_X1 U_g10465C (.ZN(g10465C),.A(I15986C));
INV_X1 U_g1980C (.ZN(g1980C),.A(g646C));
INV_X1 U_g8164C (.ZN(g8164C),.A(g2216C));
INV_X1 U_g8233C (.ZN(g8233C),.A(g2216C));
INV_X1 U_I6220C (.ZN(I6220C),.A(g883C));
INV_X1 U_I4891C (.ZN(I4891C),.A(g582C));
INV_X1 U_I4859C (.ZN(I4859C),.A(g578C));
INV_X1 U_g4212C (.ZN(g4212C),.A(I5044C));
INV_X1 U_I9479C (.ZN(I9479C),.A(g29C));
INV_X1 U_g2297C (.ZN(g2297C),.A(g865C));
INV_X1 U_g7622C (.ZN(g7622C),.A(g7067C));
INV_X1 U_I13400C (.ZN(I13400C),.A(g8236C));
INV_X1 U_g2338C (.ZN(g2338C),.A(g1909C));
INV_X1 U_g7446C (.ZN(g7446C),.A(FE_OFN86_g2176C));
INV_X1 U_g3475C (.ZN(g3475C),.A(g3056C));
INV_X1 U_g4822C (.ZN(g4822C),.A(g3706C));
INV_X1 U_g10437C (.ZN(g10437C),.A(g10333C));
INV_X1 U_g3039C (.ZN(g3039C),.A(g2310C));
INV_X1 U_I6240C (.ZN(I6240C),.A(g878C));
INV_X1 U_I9810C (.ZN(I9810C),.A(g5576C));
INV_X1 U_g2449C (.ZN(g2449C),.A(g790C));
INV_X1 U_I4783C (.ZN(I4783C),.A(g873C));
INV_X1 U_g2604C (.ZN(g2604C),.A(I5525C));
INV_X1 U_I5399C (.ZN(I5399C),.A(g895C));
INV_X1 U_g6165C (.ZN(g6165C),.A(FE_OFN100_g4421C));
INV_X1 U_I5510C (.ZN(I5510C),.A(g588C));
INV_X1 U_I5245C (.ZN(I5245C),.A(g925C));
INV_X1 U_g9505C (.ZN(g9505C),.A(FE_OFN56_g9052C));
INV_X1 U_g2268C (.ZN(g2268C),.A(g654C));
INV_X1 U_g4192C (.ZN(g4192C),.A(I5388C));
INV_X1 U_g3546C (.ZN(g3546C),.A(FE_OFN352_g109C));
INV_X4 U_g9474C (.ZN(g9474C),.A(g9331C));
INV_X1 U_g5222C (.ZN(g5222C),.A(FE_OFN153_g4640C));
INV_X1 U_g2070C (.ZN(g2070C),.A(g213C));
INV_X1 U_g3906C (.ZN(g3906C),.A(FE_OFN364_g3015C));
INV_X1 U_I4866C (.ZN(I4866C),.A(g579C));
INV_X1 U_g6256C (.ZN(g6256C),.A(g2216C));
INV_X1 U_g4176C (.ZN(g4176C),.A(g1989C));
INV_X1 U_g2331C (.ZN(g2331C),.A(g658C));
INV_X1 U_g2406C (.ZN(g2406C),.A(g1365C));
INV_X1 U_I13332C (.ZN(I13332C),.A(g8206C));
INV_X1 U_g6263C (.ZN(g6263C),.A(I9290C));
INV_X1 U_g11239C (.ZN(g11239C),.A(FE_OFN13_g10702C));
INV_X1 U_g2087C (.ZN(g2087C),.A(g225C));
INV_X1 U_g2801C (.ZN(g2801C),.A(g2117C));
INV_X1 U_g3738C (.ZN(g3738C),.A(g3062C));
INV_X1 U_g7512C (.ZN(g7512C),.A(FE_OFN86_g2176C));
INV_X1 U_g9760C (.ZN(g9760C),.A(FE_OFN33_g9454C));
INV_X1 U_g6257C (.ZN(g6257C),.A(g2169C));
INV_X1 U_g4177C (.ZN(g4177C),.A(g1990C));
INV_X1 U_g4206C (.ZN(g4206C),.A(I5579C));
INV_X1 U_g2045C (.ZN(g2045C),.A(g1811C));
INV_X1 U_g8331C (.ZN(g8331C),.A(I13373C));
INV_X1 U_I9276C (.ZN(I9276C),.A(g83C));
INV_X1 U_g8105C (.ZN(g8105C),.A(g7992C));
INV_X1 U_g2169C (.ZN(g2169C),.A(g42C));
INV_X1 U_I5395C (.ZN(I5395C),.A(g892C));
INV_X1 U_g2369C (.ZN(g2369C),.A(g617C));
INV_X1 U_g2602C (.ZN(g2602C),.A(I5497C));
INV_X1 U_g4199C (.ZN(g4199C),.A(I5418C));
INV_X1 U_g2407C (.ZN(g2407C),.A(g197C));
INV_X1 U_g9451C (.ZN(g9451C),.A(I14642C));
INV_X1 U_g5836C (.ZN(g5836C),.A(FE_OFN273_g85C));
INV_X1 U_g4207C (.ZN(g4207C),.A(I5584C));
INV_X1 U_g11083C (.ZN(g11083C),.A(g10788C));
INV_X1 U_g11348C (.ZN(g11348C),.A(g11276C));
INV_X1 U_I5815C (.ZN(I5815C),.A(g794C));
INV_X1 U_g9508C (.ZN(g9508C),.A(g9271C));
INV_X1 U_g2203C (.ZN(g2203C),.A(g677C));
INV_X1 U_g7686C (.ZN(g7686C),.A(FE_OFN85_g2176C));
INV_X1 U_I5497C (.ZN(I5497C),.A(g587C));
INV_X1 U_I13421C (.ZN(I13421C),.A(g8200C));
INV_X1 U_g4215C (.ZN(g4215C),.A(I5060C));
INV_X1 U_g6863C (.ZN(g6863C),.A(g6740C));
INV_X1 U_g2216C (.ZN(g2216C),.A(g41C));
INV_X1 U_g2028C (.ZN(g2028C),.A(g1703C));
INV_X1 U_g4336C (.ZN(g4336C),.A(g4130C));
INV_X1 U_g2564C (.ZN(g2564C),.A(g1814C));
INV_X1 U_g3705C (.ZN(g3705C),.A(FE_OFN308_I6424C));
INV_X1 U_g4065C (.ZN(g4065C),.A(g2794C));
INV_X1 U_g4887C (.ZN(g4887C),.A(I5057C));
INV_X1 U_g2609C (.ZN(g2609C),.A(I4900C));
INV_X1 U_g4934C (.ZN(g4934C),.A(g4243C));
INV_X1 U_g3814C (.ZN(g3814C),.A(g2355C));
INV_X1 U_g8564C (.ZN(g8564C),.A(I7840C));
INV_X1 U_g2571C (.ZN(g2571C),.A(g1822C));
INV_X1 U_g4195C (.ZN(g4195C),.A(I5406C));
INV_X1 U_g1975C (.ZN(g1975C),.A(g622C));
INV_X1 U_g2774C (.ZN(g2774C),.A(FE_OFN225_g2276C));
INV_X1 U_g3967C (.ZN(g3967C),.A(g3247C));
INV_X1 U_I4935C (.ZN(I4935C),.A(g585C));
INV_X1 U_g2396C (.ZN(g2396C),.A(g1389C));
INV_X1 U_g1984C (.ZN(g1984C),.A(g758C));
INV_X1 U_g11539C (.ZN(g11539C),.A(g11519C));
INV_X1 U_g2018C (.ZN(g2018C),.A(g1336C));
INV_X1 U_g2067C (.ZN(g2067C),.A(g108C));
INV_X1 U_I14323C (.ZN(I14323C),.A(g8817C));
INV_X1 U_I14299C (.ZN(I14299C),.A(g8810C));
INV_X1 U_I6277C (.ZN(I6277C),.A(g1206C));
INV_X1 U_I9237C (.ZN(I9237C),.A(g31C));
INV_X1 U_g2381C (.ZN(g2381C),.A(g1368C));
INV_X1 U_g9432C (.ZN(g9432C),.A(g9313C));
INV_X1 U_g8509C (.ZN(g8509C),.A(g8366C));
INV_X1 U_g7905C (.ZN(g7905C),.A(g7450C));
INV_X1 U_g2421C (.ZN(g2421C),.A(g1374C));
INV_X1 U_g4001C (.ZN(g4001C),.A(g3200C));
INV_X1 U_g11515C (.ZN(g11515C),.A(g11490C));
INV_X1 U_g3485C (.ZN(g3485C),.A(g1104C));
INV_X1 U_g2562C (.ZN(g2562C),.A(g1383C));
INV_X1 U_g6697C (.ZN(g6697C),.A(g4807C));
INV_X1 U_g8700C (.ZN(g8700C),.A(g8574C));
INV_X1 U_g2605C (.ZN(g2605C),.A(I4866C));
INV_X1 U_g11206C (.ZN(g11206C),.A(g10629C));
INV_X1 U_I5427C (.ZN(I5427C),.A(g913C));
INV_X1 U_I9769C (.ZN(I9769C),.A(g5287C));
INV_X1 U_g11107C (.ZN(g11107C),.A(FE_OFN7_g10702C));
INV_X1 U_I11360C (.ZN(I11360C),.A(g6351C));
INV_X1 U_g8562C (.ZN(g8562C),.A(I7825C));
INV_X1 U_g9778C (.ZN(g9778C),.A(FE_OFN63_g9474C));
INV_X1 U_g3765C (.ZN(g3765C),.A(g3120C));
INV_X1 U_g4198C (.ZN(g4198C),.A(I5414C));
INV_X1 U_I14330C (.ZN(I14330C),.A(g8819C));
INV_X1 U_g9526C (.ZN(g9526C),.A(g9256C));
INV_X1 U_I15962C (.ZN(I15962C),.A(g10405C));
INV_X1 U_g3069C (.ZN(g3069C),.A(I6277C));
INV_X1 U_I15500C (.ZN(I15500C),.A(g10019C));
INV_X1 U_I5047C (.ZN(I5047C),.A(g1185C));
INV_X1 U_g2074C (.ZN(g2074C),.A(g1377C));
INV_X1 U_I16507C (.ZN(I16507C),.A(g10712C));
INV_X1 U_g6942C (.ZN(g6942C),.A(I7840C));
INV_X1 U_g4211C (.ZN(g4211C),.A(I5041C));
INV_X1 U_g6432C (.ZN(g6432C),.A(FE_OFN219_g5557C));
INV_X1 U_g7908C (.ZN(g7908C),.A(g7454C));
INV_X1 U_g9764C (.ZN(g9764C),.A(FE_OFN59_g9432C));
INV_X1 U_g3291C (.ZN(g3291C),.A(g2161C));
INV_X1 U_g3207C (.ZN(g3207C),.A(g2439C));
INV_X1 U_g2126C (.ZN(g2126C),.A(g12C));
INV_X1 U_I15514C (.ZN(I15514C),.A(g10007C));
INV_X1 U_I15507C (.ZN(I15507C),.A(g10001C));
INV_X1 U_g1964C (.ZN(g1964C),.A(g114C));
INV_X1 U_g10387C (.ZN(g10387C),.A(g10357C));
INV_X1 U_g11163C (.ZN(g11163C),.A(I16717C));
INV_X1 U_g8688C (.ZN(g8688C),.A(g8507C));
INV_X1 U_g8976C (.ZN(g8976C),.A(I14323C));
INV_X1 U_g2608C (.ZN(g2608C),.A(I4891C));
INV_X1 U_g7450C (.ZN(g7450C),.A(FE_OFN87_g2176C));
INV_X1 U_g4200C (.ZN(g4200C),.A(I5424C));
INV_X1 U_g2023C (.ZN(g2023C),.A(g1357C));
INV_X1 U_g7379C (.ZN(g7379C),.A(g6863C));
INV_X1 U_I13427C (.ZN(I13427C),.A(g8241C));
INV_X1 U_I7752C (.ZN(I7752C),.A(g3407C));
INV_X1 U_g4191C (.ZN(g4191C),.A(I5383C));
INV_X1 U_g1989C (.ZN(g1989C),.A(g770C));
INV_X1 U_g3408C (.ZN(g3408C),.A(g3108C));
INV_X1 U_g2451C (.ZN(g2451C),.A(g248C));
INV_X1 U_g8220C (.ZN(g8220C),.A(FE_OFN199_g7697C));
INV_X1 U_g3943C (.ZN(g3943C),.A(g627C));
INV_X1 U_I14295C (.ZN(I14295C),.A(g8806C));
INV_X1 U_g7981C (.ZN(g7981C),.A(g7624C));
INV_X1 U_g6949C (.ZN(g6949C),.A(I7847C));
INV_X1 U_g8977C (.ZN(g8977C),.A(I14295C));
INV_X1 U_g9082C (.ZN(g9082C),.A(FE_OFN76_g8700C));
INV_X1 U_g4811C (.ZN(g4811C),.A(g3661C));
INV_X1 U_g10379C (.ZN(g10379C),.A(I15861C));
INV_X1 U_g7680C (.ZN(g7680C),.A(FE_OFN87_g2176C));
INV_X1 U_g8327C (.ZN(g8327C),.A(g8164C));
INV_X1 U_I13385C (.ZN(I13385C),.A(g8230C));
INV_X1 U_g7744C (.ZN(g7744C),.A(g1962C));
INV_X1 U_g8146C (.ZN(g8146C),.A(FE_OFN330_g7638C));
INV_X1 U_I5057C (.ZN(I5057C),.A(g1961C));
INV_X1 U_I8503C (.ZN(I8503C),.A(FE_OFN184_I7048C));
INV_X1 U_g2034C (.ZN(g2034C),.A(g1766C));
INV_X1 U_g8103C (.ZN(g8103C),.A(g7994C));
INV_X1 U_g2434C (.ZN(g2434C),.A(g1362C));
INV_X1 U_g3913C (.ZN(g3913C),.A(g3121C));
INV_X1 U_g6702C (.ZN(g6702C),.A(FE_OFN117_g4807C));
INV_X1 U_g4880C (.ZN(g4880C),.A(FE_OFN292_g3015C));
INV_X1 U_g8696C (.ZN(g8696C),.A(g8488C));
INV_X1 U_I14309C (.ZN(I14309C),.A(g8813C));
INV_X1 U_g2347C (.ZN(g2347C),.A(g1945C));
INV_X1 U_g6276C (.ZN(g6276C),.A(I9329C));
INV_X1 U_g4243C (.ZN(g4243C),.A(g3524C));
INV_X1 U_I9259C (.ZN(I9259C),.A(g89C));
INV_X1 U_g7574C (.ZN(g7574C),.A(FE_OFN80_g2175C));
INV_X1 U_g8316C (.ZN(g8316C),.A(I13332C));
INV_X1 U_g8565C (.ZN(g8565C),.A(I7847C));
INV_X1 U_g8347C (.ZN(g8347C),.A(I13421C));
INV_X1 U_g1962C (.ZN(g1962C),.A(g27C));
INV_X1 U_g2601C (.ZN(g2601C),.A(I4859C));
INV_X1 U_g4213C (.ZN(g4213C),.A(I5047C));
INV_X1 U_g6277C (.ZN(g6277C),.A(I9349C));
INV_X1 U_g2060C (.ZN(g2060C),.A(g1380C));
INV_X1 U_g6617C (.ZN(g6617C),.A(g6019C));
INV_X1 U_I13338C (.ZN(I13338C),.A(g8210C));
INV_X1 U_I15861C (.ZN(I15861C),.A(g10339C));
INV_X1 U_I5525C (.ZN(I5525C),.A(g589C));
INV_X1 U_g4456C (.ZN(g4456C),.A(FE_OFN234_g2024C));
INV_X1 U_g2479C (.ZN(g2479C),.A(g26C));
INV_X1 U_I16220C (.ZN(I16220C),.A(g10502C));
INV_X1 U_g9814C (.ZN(g9814C),.A(FE_OFN70_g9490C));
INV_X1 U_g3068C (.ZN(g3068C),.A(g2303C));
INV_X1 U_g9773C (.ZN(g9773C),.A(g9474C));
INV_X1 U_g5200C (.ZN(g5200C),.A(g4567C));
INV_X1 U_g4457C (.ZN(g4457C),.A(FE_OFN137_g3829C));
INV_X1 U_g4193C (.ZN(g4193C),.A(I5395C));
INV_X1 U_g10461C (.ZN(g10461C),.A(I15974C));
INV_X1 U_I5020C (.ZN(I5020C),.A(g1176C));
INV_X1 U_g1969C (.ZN(g1969C),.A(g456C));
INV_X1 U_I9293C (.ZN(I9293C),.A(g92C));
INV_X1 U_I9329C (.ZN(I9329C),.A(g94C));
INV_X1 U_g7903C (.ZN(g7903C),.A(g7446C));
INV_X1 U_I9221C (.ZN(I9221C),.A(g30C));
INV_X1 U_g4525C (.ZN(g4525C),.A(FE_OFN229_g3880C));
INV_X1 U_g2475C (.ZN(g2475C),.A(g192C));
INV_X1 U_g1988C (.ZN(g1988C),.A(g766C));
INV_X1 U_g11203C (.ZN(g11203C),.A(FE_OFN20_g10702C));
INV_X1 U_g4158C (.ZN(g4158C),.A(g3304C));
INV_X1 U_g6557C (.ZN(g6557C),.A(FE_OFN217_g5013C));
INV_X1 U_g2603C (.ZN(g2603C),.A(I5510C));
INV_X1 U_I5410C (.ZN(I5410C),.A(g901C));
INV_X1 U_g10459C (.ZN(g10459C),.A(I15968C));
INV_X1 U_I9349C (.ZN(I9349C),.A(g95C));
INV_X1 U_g6955C (.ZN(g6955C),.A(I7852C));
INV_X1 U_I15290C (.ZN(I15290C),.A(g9974C));
INV_X1 U_g6254C (.ZN(g6254C),.A(I9221C));
INV_X1 U_g4174C (.ZN(g4174C),.A(g1987C));
INV_X1 U_g10444C (.ZN(g10444C),.A(g10325C));
INV_X1 U_I14642C (.ZN(I14642C),.A(g9088C));
INV_X1 U_g4180C (.ZN(g4180C),.A(g1993C));
INV_X1 U_g7917C (.ZN(g7917C),.A(g7497C));
INV_X1 U_g2986C (.ZN(g2986C),.A(I6220C));
INV_X1 U_g9473C (.ZN(g9473C),.A(g9082C));
INV_X1 U_g1965C (.ZN(g1965C),.A(g119C));
INV_X1 U_g11547C (.ZN(g11547C),.A(FE_OFN27_g11519C));
INV_X1 U_g2503C (.ZN(g2503C),.A(g1872C));
INV_X1 U_I9352C (.ZN(I9352C),.A(g28C));
INV_X1 U_I9717C (.ZN(I9717C),.A(FE_OFN97_I8869C));
INV_X1 U_g2224C (.ZN(g2224C),.A(g695C));
INV_X1 U_g7454C (.ZN(g7454C),.A(g2176C));
INV_X1 U_g4204C (.ZN(g4204C),.A(I5445C));
INV_X1 U_g8561C (.ZN(g8561C),.A(I7817C));
INV_X1 U_g8986C (.ZN(g8986C),.A(I14330C));
INV_X1 U_I15956C (.ZN(I15956C),.A(g10402C));
INV_X1 U_I15980C (.ZN(I15980C),.A(g10414C));
AND2_X1 U_g11103C (.ZN(g11103C),.A2(g10937C),.A1(g2250C));
AND2_X1 U_g9900C (.ZN(g9900C),.A2(g8327C),.A1(g9088C));
AND2_X1 U_g11095C (.ZN(g11095C),.A2(FE_OFN4_g10950C),.A1(g845C));
AND2_X2 U_g3880C (.ZN(g3880C),.A2(g2023C),.A1(FE_OFN235_g2024C));
AND2_X1 U_g4973C (.ZN(g4973C),.A2(g4467C),.A1(g1645C));
AND2_X1 U_g7389C (.ZN(g7389C),.A2(FE_OFN226_g3880C),.A1(g5852C));
AND2_X1 U_g7888C (.ZN(g7888C),.A2(FE_OFN334_g7045C),.A1(g7465C));
AND2_X1 U_g4969C (.ZN(g4969C),.A2(g4457C),.A1(g1642C));
AND2_X1 U_g8224C (.ZN(g8224C),.A2(g7949C),.A1(g1882C));
AND2_X1 U_g2892C (.ZN(g2892C),.A2(g1976C),.A1(g1980C));
AND2_X1 U_g5686C (.ZN(g5686C),.A2(FE_OFN365_g5361C),.A1(g158C));
AND2_X1 U_g10308C (.ZN(g10308C),.A2(g9082C),.A1(g10013C));
AND2_X1 U_g4123C (.ZN(g4123C),.A2(g2424C),.A1(g1781C));
AND2_X1 U_g8120C (.ZN(g8120C),.A2(g7949C),.A1(g1909C));
AND2_X1 U_g6788C (.ZN(g6788C),.A2(FE_OFN320_g5361C),.A1(g287C));
AND2_X1 U_g5598C (.ZN(g5598C),.A2(g4824C),.A1(g778C));
AND2_X1 U_g9694C (.ZN(g9694C),.A2(FE_OFN59_g9432C),.A1(g278C));
AND2_X1 U_g10495C (.ZN(g10495C),.A2(FE_OFN234_g2024C),.A1(g10431C));
AND2_X1 U_g2945C (.ZN(g2945C),.A2(g1684C),.A1(FE_OFN241_g1690C));
AND2_X1 U_g11190C (.ZN(g11190C),.A2(g10927C),.A1(g4752C));
AND2_X1 U_g8789C (.ZN(g8789C),.A2(FE_OFN331_g8696C),.A1(g8639C));
AND2_X1 U_g9852C (.ZN(g9852C),.A2(g9563C),.A1(g9728C));
AND2_X1 U_g5625C (.ZN(g5625C),.A2(g5627C),.A1(g1053C));
AND2_X1 U_g4875C (.ZN(g4875C),.A2(g4673C),.A1(g995C));
AND2_X1 U_g9701C (.ZN(g9701C),.A2(g9474C),.A1(g1574C));
AND2_X1 U_g7138C (.ZN(g7138C),.A2(g6718C),.A1(g5201C));
AND2_X1 U_g10752C (.ZN(g10752C),.A2(FE_OFN103_g3586C),.A1(g10599C));
AND2_X1 U_g11211C (.ZN(g11211C),.A2(g5503C),.A1(g11058C));
AND2_X1 U_g11024C (.ZN(g11024C),.A2(g10702C),.A1(g435C));
AND2_X1 U_g8547C (.ZN(g8547C),.A2(FE_OFN211_g7246C),.A1(g8307C));
AND2_X1 U_g10669C (.ZN(g10669C),.A2(g9473C),.A1(g10408C));
AND2_X1 U_g7707C (.ZN(g7707C),.A2(FE_OFN191_g6488C),.A1(g691C));
AND2_X1 U_g4884C (.ZN(g4884C),.A2(g1845C),.A1(g3813C));
AND2_X1 U_g4839C (.ZN(g4839C),.A2(g2355C),.A1(g225C));
AND2_X1 U_g9870C (.ZN(g9870C),.A2(g9802C),.A1(g1561C));
AND2_X1 U_g6640C (.ZN(g6640C),.A2(g5808C),.A1(g86C));
AND2_X1 U_g9650C (.ZN(g9650C),.A2(FE_OFN40_g9240C),.A1(g986C));
AND2_X1 U_g5687C (.ZN(g5687C),.A2(FE_OFN365_g5361C),.A1(g139C));
AND2_X1 U_g7957C (.ZN(g7957C),.A2(g7527C),.A1(g79C));
AND2_X1 U_g3512C (.ZN(g3512C),.A2(g1845C),.A1(g2050C));
AND2_X1 U_g8244C (.ZN(g8244C),.A2(FE_OFN310_g4336C),.A1(g7054C));
AND2_X1 U_g7449C (.ZN(g7449C),.A2(FE_OFN221_g3440C),.A1(g6548C));
AND2_X1 U_g4235C (.ZN(g4235C),.A2(FE_OFN347_g3914C),.A1(g1011C));
AND2_X1 U_g4343C (.ZN(g4343C),.A2(FE_OFN287_g3586C),.A1(g345C));
AND2_X1 U_g11296C (.ZN(g11296C),.A2(g11239C),.A1(g4561C));
AND2_X1 U_g9594C (.ZN(g9594C),.A2(g9292C),.A1(g1C));
AND2_X1 U_g6829C (.ZN(g6829C),.A2(FE_OFN179_g5354C),.A1(g213C));
AND2_X1 U_g4334C (.ZN(g4334C),.A2(FE_OFN351_g3913C),.A1(g1160C));
AND2_X1 U_g9943C (.ZN(g9943C),.A2(FE_OFN67_g9367C),.A1(g9923C));
AND2_X1 U_g5525C (.ZN(g5525C),.A2(g4292C),.A1(g1721C));
AND2_X1 U_g4548C (.ZN(g4548C),.A2(g4002C),.A1(g440C));
AND3_X1 U_g8876C (.ZN(g8876C),.A3(FE_OFN73_g8858C),.A2(FE_OFN93_g2216C),.A1(g8105C));
AND2_X1 U_g6733C (.ZN(g6733C),.A2(FE_OFN322_g4449C),.A1(g4488C));
AND2_X1 U_g4804C (.ZN(g4804C),.A2(g4010C),.A1(g476C));
AND2_X1 U_g10705C (.ZN(g10705C),.A2(FE_OFN131_g3015C),.A1(g10564C));
AND2_X1 U_g9934C (.ZN(g9934C),.A2(g9624C),.A1(g9913C));
AND2_X1 U_g6225C (.ZN(g6225C),.A2(g5613C),.A1(g566C));
AND2_X1 U_g6324C (.ZN(g6324C),.A2(FE_OFN116_g4807C),.A1(g1240C));
AND2_X1 U_g10686C (.ZN(g10686C),.A2(FE_OFN136_g3863C),.A1(g10385C));
AND2_X1 U_g6540C (.ZN(g6540C),.A2(g6081C),.A1(g1223C));
AND2_X1 U_g8663C (.ZN(g8663C),.A2(FE_OFN292_g3015C),.A1(g8270C));
AND2_X1 U_g11581C (.ZN(g11581C),.A2(g11539C),.A1(g1308C));
AND2_X1 U_g6206C (.ZN(g6206C),.A2(g5613C),.A1(g560C));
AND2_X1 U_g4518C (.ZN(g4518C),.A2(g4002C),.A1(g452C));
AND2_X1 U_g3989C (.ZN(g3989C),.A2(FE_OFN359_g18C),.A1(g248C));
AND2_X1 U_g7730C (.ZN(g7730C),.A2(g2347C),.A1(g7260C));
AND2_X1 U_g5174C (.ZN(g5174C),.A2(FE_OFN303_g4678C),.A1(g1235C));
AND2_X1 U_g7504C (.ZN(g7504C),.A2(g67C),.A1(FE_OFN86_g2176C));
AND2_X1 U_g7185C (.ZN(g7185C),.A2(FE_OFN213_g6003C),.A1(g1887C));
AND2_X1 U_g2563C (.ZN(g2563C),.A2(I5690C),.A1(I5689C));
AND2_X1 U_g7881C (.ZN(g7881C),.A2(FE_OFN366_g3521C),.A1(g5295C));
AND2_X1 U_g11070C (.ZN(g11070C),.A2(g10788C),.A1(g2008C));
AND2_X1 U_g9859C (.ZN(g9859C),.A2(g9579C),.A1(g9736C));
AND3_X1 U_g8877C (.ZN(g8877C),.A3(FE_OFN73_g8858C),.A2(FE_OFN92_g2216C),.A1(g8103C));
AND2_X1 U_g11590C (.ZN(g11590C),.A2(g11561C),.A1(g2274C));
AND2_X1 U_g6199C (.ZN(g6199C),.A2(FE_OFN289_g4679C),.A1(g557C));
AND2_X1 U_g9266C (.ZN(g9266C),.A2(FE_OFN325_g18C),.A1(g8932C));
AND2_X1 U_g5545C (.ZN(g5545C),.A2(g4292C),.A1(g1730C));
AND2_X1 U_g5180C (.ZN(g5180C),.A2(g810C),.A1(g814C));
AND2_X1 U_g5591C (.ZN(g5591C),.A2(FE_OFN367_g3521C),.A1(g1615C));
AND2_X1 U_g8556C (.ZN(g8556C),.A2(FE_OFN189_g7638C),.A1(g8412C));
AND2_X1 U_g11094C (.ZN(g11094C),.A2(g10883C),.A1(g374C));
AND2_X1 U_g5853C (.ZN(g5853C),.A2(g1927C),.A1(g5044C));
AND2_X1 U_g6245C (.ZN(g6245C),.A2(FE_OFN289_g4679C),.A1(g575C));
AND2_X1 U_g4360C (.ZN(g4360C),.A2(g3523C),.A1(g1861C));
AND3_X1 U_g8930C (.ZN(g8930C),.A3(g8828C),.A2(FE_OFN95_g2216C),.A1(g8100C));
AND2_X1 U_g5507C (.ZN(g5507C),.A2(FE_OFN357_g3521C),.A1(g563C));
AND2_X1 U_g11150C (.ZN(g11150C),.A2(g10788C),.A1(g3087C));
AND2_X1 U_g8464C (.ZN(g8464C),.A2(FE_OFN210_g7246C),.A1(g8302C));
AND2_X1 U_g9692C (.ZN(g9692C),.A2(FE_OFN59_g9432C),.A1(g272C));
AND2_X1 U_g4996C (.ZN(g4996C),.A2(FE_OFN146_g4682C),.A1(g1428C));
AND2_X1 U_g7131C (.ZN(g7131C),.A2(g6702C),.A1(g5174C));
AND2_X1 U_g11019C (.ZN(g11019C),.A2(FE_OFN7_g10702C),.A1(g421C));
AND2_X1 U_g9960C (.ZN(g9960C),.A2(FE_OFN280_g9536C),.A1(g9951C));
AND2_X1 U_g11196C (.ZN(g11196C),.A2(FE_OFN15_g10702C),.A1(g4770C));
AND2_X1 U_g11018C (.ZN(g11018C),.A2(FE_OFN7_g10702C),.A1(g6485C));
AND2_X1 U_g6819C (.ZN(g6819C),.A2(FE_OFN179_g5354C),.A1(g243C));
AND2_X1 U_g10595C (.ZN(g10595C),.A2(FE_OFN369_g4525C),.A1(g10550C));
AND2_X1 U_g10494C (.ZN(g10494C),.A2(g2024C),.A1(g10433C));
AND2_X1 U_g10623C (.ZN(g10623C),.A2(FE_OFN370_g4525C),.A1(g10544C));
AND2_X1 U_g4878C (.ZN(g4878C),.A2(g3523C),.A1(g1868C));
AND2_X1 U_g5204C (.ZN(g5204C),.A2(g2126C),.A1(g4838C));
AND2_X1 U_g8844C (.ZN(g8844C),.A2(g8709C),.A1(g8609C));
AND2_X1 U_g6701C (.ZN(g6701C),.A2(g4381C),.A1(g6185C));
AND2_X1 U_g10782C (.ZN(g10782C),.A2(g4467C),.A1(g10725C));
AND2_X1 U_g5100C (.ZN(g5100C),.A2(g4608C),.A1(g1791C));
AND2_X1 U_g4882C (.ZN(g4882C),.A2(FE_OFN293_g3015C),.A1(g1089C));
AND2_X1 U_g8731C (.ZN(g8731C),.A2(g7918C),.A1(g8236C));
AND2_X1 U_g6215C (.ZN(g6215C),.A2(g5128C),.A1(g1504C));
AND2_X1 U_g6886C (.ZN(g6886C),.A2(FE_OFN213_g6003C),.A1(g1932C));
AND2_X4 U_g3586C (.ZN(g3586C),.A2(I6260C),.A1(g1703C));
AND2_X1 U_g8557C (.ZN(g8557C),.A2(g7638C),.A1(g8415C));
AND3_X1 U_g8966C (.ZN(g8966C),.A3(g8849C),.A2(FE_OFN93_g2216C),.A1(g8081C));
AND2_X1 U_g8071C (.ZN(g8071C),.A2(FE_OFN199_g7697C),.A1(g691C));
AND2_X1 U_g11597C (.ZN(g11597C),.A2(FE_OFN99_g4421C),.A1(g11549C));
AND2_X1 U_g9828C (.ZN(g9828C),.A2(g9785C),.A1(g9722C));
AND2_X1 U_g2918C (.ZN(g2918C),.A2(g1672C),.A1(FE_OFN241_g1690C));
AND2_X1 U_g9830C (.ZN(g9830C),.A2(FE_OFN34_g9785C),.A1(g9725C));
AND3_X1 U_g8955C (.ZN(g8955C),.A3(g8828C),.A2(FE_OFN95_g2216C),.A1(g8110C));
AND2_X1 U_g9592C (.ZN(g9592C),.A2(g9292C),.A1(g4C));
AND2_X1 U_g5123C (.ZN(g5123C),.A2(g3906C),.A1(g1618C));
AND2_X1 U_g7059C (.ZN(g7059C),.A2(g6354C),.A1(g6078C));
AND2_X1 U_g8254C (.ZN(g8254C),.A2(g7907C),.A1(g936C));
AND2_X1 U_g7459C (.ZN(g7459C),.A2(g55C),.A1(FE_OFN86_g2176C));
AND2_X1 U_g11102C (.ZN(g11102C),.A2(FE_OFN3_g10950C),.A1(g861C));
AND2_X1 U_g7718C (.ZN(g7718C),.A2(FE_OFN191_g6488C),.A1(g709C));
AND2_X1 U_g7535C (.ZN(g7535C),.A2(g49C),.A1(FE_OFN86_g2176C));
AND2_X1 U_g9703C (.ZN(g9703C),.A2(g9474C),.A1(g1577C));
AND2_X1 U_g5528C (.ZN(g5528C),.A2(FE_OFN357_g3521C),.A1(g569C));
AND2_X1 U_g9932C (.ZN(g9932C),.A2(g9624C),.A1(g9911C));
AND2_X1 U_g5530C (.ZN(g5530C),.A2(FE_OFN290_g4880C),.A1(g1636C));
AND2_X1 U_g3506C (.ZN(g3506C),.A2(g2760C),.A1(g986C));
AND2_X1 U_g8769C (.ZN(g8769C),.A2(FE_OFN304_g5151C),.A1(g8629C));
AND2_X1 U_g6887C (.ZN(g6887C),.A2(g6557C),.A1(g6187C));
AND2_X1 U_g6228C (.ZN(g6228C),.A2(g713C),.A1(g5605C));
AND2_X1 U_g6322C (.ZN(g6322C),.A2(FE_OFN116_g4807C),.A1(g1275C));
AND2_X1 U_g3111C (.ZN(g3111C),.A2(I6338C),.A1(I6337C));
AND3_X1 U_g8967C (.ZN(g8967C),.A3(g8849C),.A2(FE_OFN281_g2216C),.A1(g8085C));
AND2_X1 U_g5010C (.ZN(g5010C),.A2(FE_OFN153_g4640C),.A1(g1458C));
AND2_X1 U_g3275C (.ZN(g3275C),.A2(FE_OFN266_g18C),.A1(g115C));
AND2_X1 U_g10809C (.ZN(g10809C),.A2(g10702C),.A1(g4811C));
AND2_X1 U_g2895C (.ZN(g2895C),.A2(g1678C),.A1(FE_OFN336_g1690C));
AND2_X1 U_g7721C (.ZN(g7721C),.A2(g6488C),.A1(g736C));
AND2_X1 U_g9866C (.ZN(g9866C),.A2(g9802C),.A1(g1549C));
AND2_X1 U_g9716C (.ZN(g9716C),.A2(FE_OFN70_g9490C),.A1(g1534C));
AND2_X1 U_g10808C (.ZN(g10808C),.A2(FE_OFN137_g3829C),.A1(g10744C));
AND2_X1 U_g3374C (.ZN(g3374C),.A2(g3047C),.A1(g1231C));
AND2_X1 U_g4492C (.ZN(g4492C),.A2(g3685C),.A1(FE_OFN253_g1786C));
AND2_X1 U_g8822C (.ZN(g8822C),.A2(FE_OFN328_g8709C),.A1(g8614C));
AND2_X1 U_g10560C (.ZN(g10560C),.A2(FE_OFN369_g4525C),.A1(g10369C));
AND3_X1 U_g11456C (.ZN(g11456C),.A3(g11348C),.A2(g2801C),.A1(g3765C));
AND2_X1 U_g9848C (.ZN(g9848C),.A2(g9579C),.A1(g9724C));
AND2_X1 U_g4714C (.ZN(g4714C),.A2(g3943C),.A1(g646C));
AND2_X1 U_g6550C (.ZN(g6550C),.A2(g6081C),.A1(g1231C));
AND2_X1 U_g5172C (.ZN(g5172C),.A2(g818C),.A1(g822C));
AND2_X1 U_g10642C (.ZN(g10642C),.A2(g3829C),.A1(g10385C));
AND2_X1 U_g3284C (.ZN(g3284C),.A2(g677C),.A1(g2531C));
AND2_X1 U_g9699C (.ZN(g9699C),.A2(FE_OFN59_g9432C),.A1(g284C));
AND2_X1 U_g9855C (.ZN(g9855C),.A2(g9764C),.A1(g302C));
AND2_X1 U_g5618C (.ZN(g5618C),.A2(FE_OFN367_g3521C),.A1(g1630C));
AND2_X1 U_g6891C (.ZN(g6891C),.A2(g6003C),.A1(g1950C));
AND2_X1 U_g7940C (.ZN(g7940C),.A2(FE_OFN292_g3015C),.A1(g5319C));
AND2_X1 U_g11085C (.ZN(g11085C),.A2(g10927C),.A1(g312C));
AND2_X1 U_g4736C (.ZN(g4736C),.A2(FE_OFN300_g4002C),.A1(g396C));
AND2_X1 U_g4968C (.ZN(g4968C),.A2(FE_OFN146_g4682C),.A1(g1432C));
AND2_X1 U_g8837C (.ZN(g8837C),.A2(FE_OFN331_g8696C),.A1(g8646C));
AND2_X1 U_g9644C (.ZN(g9644C),.A2(FE_OFN45_g9125C),.A1(g1182C));
AND2_X1 U_g5804C (.ZN(g5804C),.A2(g5261C),.A1(g1546C));
AND2_X1 U_g8462C (.ZN(g8462C),.A2(FE_OFN211_g7246C),.A1(g8300C));
AND4_X1 U_I6330C (.ZN(I6330C),.A4(g2570C),.A3(g2562C),.A2(g2556C),.A1(g2549C));
AND2_X1 U_g11156C (.ZN(g11156C),.A2(FE_OFN278_g10927C),.A1(g333C));
AND2_X1 U_g6342C (.ZN(g6342C),.A2(FE_OFN319_g5361C),.A1(g293C));
AND2_X1 U_g9867C (.ZN(g9867C),.A2(g9802C),.A1(g1552C));
AND2_X1 U_g9717C (.ZN(g9717C),.A2(FE_OFN70_g9490C),.A1(g1537C));
AND2_X1 U_g4871C (.ZN(g4871C),.A2(g3523C),.A1(g1864C));
AND2_X1 U_g10454C (.ZN(g10454C),.A2(FE_OFN235_g2024C),.A1(g10435C));
AND2_X1 U_g4722C (.ZN(g4722C),.A2(FE_OFN300_g4002C),.A1(g426C));
AND2_X1 U_g7741C (.ZN(g7741C),.A2(g3880C),.A1(g5824C));
AND2_X1 U_g4500C (.ZN(g4500C),.A2(FE_OFN291_g4880C),.A1(g1357C));
AND2_X1 U_g9386C (.ZN(g9386C),.A2(FE_OFN47_g9151C),.A1(g1327C));
AND2_X1 U_g8842C (.ZN(g8842C),.A2(FE_OFN328_g8709C),.A1(g8607C));
AND2_X1 U_g9599C (.ZN(g9599C),.A2(FE_OFN71_g9292C),.A1(g8C));
AND2_X4 U_g9274C (.ZN(g9274C),.A2(FE_OFN275_g48C),.A1(g8974C));
AND2_X1 U_g5518C (.ZN(g5518C),.A2(FE_OFN357_g3521C),.A1(g566C));
AND2_X1 U_g9614C (.ZN(g9614C),.A2(FE_OFN51_g9111C),.A1(g1197C));
AND2_X1 U_g4838C (.ZN(g4838C),.A2(g4122C),.A1(g3275C));
AND2_X4 U_g9125C (.ZN(g9125C),.A2(FE_OFN276_g48C),.A1(g8966C));
AND2_X1 U_g7217C (.ZN(g7217C),.A2(g6432C),.A1(g4610C));
AND2_X1 U_g11557C (.ZN(g11557C),.A2(g11519C),.A1(g1791C));
AND2_X1 U_g2911C (.ZN(g2911C),.A2(g1675C),.A1(FE_OFN336_g1690C));
AND2_X1 U_g11210C (.ZN(g11210C),.A2(FE_OFN204_g3664C),.A1(g10886C));
AND2_X1 U_g7466C (.ZN(g7466C),.A2(g58C),.A1(g2176C));
AND2_X1 U_g9939C (.ZN(g9939C),.A2(FE_OFN67_g9367C),.A1(g9918C));
AND2_X1 U_g11279C (.ZN(g11279C),.A2(g11203C),.A1(g4784C));
AND3_X1 U_g10518C (.ZN(g10518C),.A3(I16145C),.A2(g10440C),.A1(g10513C));
AND2_X1 U_g4477C (.ZN(g4477C),.A2(g3913C),.A1(g1129C));
AND2_X1 U_g7055C (.ZN(g7055C),.A2(g6586C),.A1(g5004C));
AND2_X1 U_g5264C (.ZN(g5264C),.A2(g4776C),.A1(g1095C));
AND2_X1 U_g6329C (.ZN(g6329C),.A2(FE_OFN115_g4807C),.A1(g1265C));
AND2_X1 U_g6828C (.ZN(g6828C),.A2(FE_OFN179_g5354C),.A1(g1377C));
AND2_X1 U_g8176C (.ZN(g8176C),.A2(FE_OFN89_I11360C),.A1(g40C));
AND2_X1 U_g6830C (.ZN(g6830C),.A2(FE_OFN179_g5354C),.A1(g1380C));
AND2_X1 U_g8005C (.ZN(g8005C),.A2(FE_OFN334_g7045C),.A1(g7510C));
AND2_X1 U_g4099C (.ZN(g4099C),.A2(g3281C),.A1(g770C));
AND2_X1 U_g11601C (.ZN(g11601C),.A2(g11575C),.A1(g1351C));
AND2_X1 U_g11187C (.ZN(g11187C),.A2(FE_OFN10_g10702C),.A1(g4727C));
AND2_X1 U_g6746C (.ZN(g6746C),.A2(FE_OFN218_g5557C),.A1(g6228C));
AND2_X1 U_g6221C (.ZN(g6221C),.A2(g5598C),.A1(g782C));
AND2_X1 U_g8765C (.ZN(g8765C),.A2(FE_OFN304_g5151C),.A1(g8630C));
AND2_X1 U_g9622C (.ZN(g9622C),.A2(FE_OFN51_g9111C),.A1(g1200C));
AND2_X1 U_g11143C (.ZN(g11143C),.A2(g4567C),.A1(g10923C));
AND2_X1 U_g9904C (.ZN(g9904C),.A2(g9676C),.A1(g9886C));
AND2_X1 U_g8733C (.ZN(g8733C),.A2(g7920C),.A1(g8241C));
AND3_X1 U_g8974C (.ZN(g8974C),.A3(FE_OFN73_g8858C),.A2(FE_OFN93_g2216C),.A1(g8094C));
AND2_X1 U_g6624C (.ZN(g6624C),.A2(FE_OFN282_g6165C),.A1(g348C));
AND2_X1 U_g11169C (.ZN(g11169C),.A2(FE_OFN8_g10702C),.A1(g530C));
AND2_X1 U_g8073C (.ZN(g8073C),.A2(FE_OFN199_g7697C),.A1(g709C));
AND2_X1 U_g9841C (.ZN(g9841C),.A2(g9512C),.A1(g9706C));
AND2_X1 U_g5882C (.ZN(g5882C),.A2(FE_OFN141_g3829C),.A1(g5592C));
AND2_X1 U_g8796C (.ZN(g8796C),.A2(FE_OFN331_g8696C),.A1(g8645C));
AND2_X1 U_g11168C (.ZN(g11168C),.A2(FE_OFN7_g10702C),.A1(g534C));
AND2_X1 U_g4269C (.ZN(g4269C),.A2(FE_OFN347_g3914C),.A1(g1015C));
AND2_X1 U_g5271C (.ZN(g5271C),.A2(FE_OFN335_g4737C),.A1(g727C));
AND2_X1 U_g10348C (.ZN(g10348C),.A2(g3705C),.A1(I15500C));
AND2_X1 U_g5611C (.ZN(g5611C),.A2(g4880C),.A1(g1047C));
AND2_X1 U_g8069C (.ZN(g8069C),.A2(FE_OFN198_g7697C),.A1(g673C));
AND2_X1 U_g9695C (.ZN(g9695C),.A2(g9474C),.A1(g1567C));
AND2_X1 U_g10304C (.ZN(g10304C),.A2(g9291C),.A1(g10001C));
AND2_X1 U_g8469C (.ZN(g8469C),.A2(FE_OFN211_g7246C),.A1(g8305C));
AND2_X1 U_g4712C (.ZN(g4712C),.A2(FE_OFN297_g3015C),.A1(g1071C));
AND2_X1 U_g6576C (.ZN(g6576C),.A2(g5503C),.A1(g5762C));
AND2_X1 U_g10622C (.ZN(g10622C),.A2(FE_OFN369_g4525C),.A1(g10496C));
AND2_X1 U_g11015C (.ZN(g11015C),.A2(FE_OFN18_g10702C),.A1(g5217C));
AND2_X1 U_g5674C (.ZN(g5674C),.A2(FE_OFN365_g5361C),.A1(g148C));
AND2_X1 U_g9359C (.ZN(g9359C),.A2(FE_OFN52_g9173C),.A1(g1308C));
AND2_X2 U_g9223C (.ZN(g9223C),.A2(g8960C),.A1(FE_OFN277_g48C));
AND2_X1 U_g11556C (.ZN(g11556C),.A2(g11519C),.A1(g1786C));
AND2_X1 U_g9858C (.ZN(g9858C),.A2(g9778C),.A1(g1595C));
AND2_X1 U_g5541C (.ZN(g5541C),.A2(g3521C),.A1(g575C));
AND2_X1 U_g4534C (.ZN(g4534C),.A2(FE_OFN344_g3586C),.A1(g363C));
AND2_X1 U_g6198C (.ZN(g6198C),.A2(g5128C),.A1(g1499C));
AND2_X1 U_g6747C (.ZN(g6747C),.A2(g5897C),.A1(g2214C));
AND2_X1 U_g6699C (.ZN(g6699C),.A2(FE_OFN111_g3914C),.A1(g6177C));
AND2_X1 U_g6855C (.ZN(g6855C),.A2(g6392C),.A1(g1964C));
AND2_X1 U_g3804C (.ZN(g3804C),.A2(g2203C),.A1(g3098C));
AND2_X1 U_g5680C (.ZN(g5680C),.A2(FE_OFN164_g5361C),.A1(g153C));
AND2_X1 U_g9642C (.ZN(g9642C),.A2(FE_OFN40_g9240C),.A1(g981C));
AND2_X1 U_g5744C (.ZN(g5744C),.A2(FE_OFN321_g5261C),.A1(g1528C));
AND2_X1 U_g10333C (.ZN(g10333C),.A2(FE_OFN267_g109C),.A1(I15500C));
AND2_X1 U_g8399C (.ZN(g8399C),.A2(g8220C),.A1(g5266C));
AND2_X1 U_g9447C (.ZN(g9447C),.A2(FE_OFN49_g9030C),.A1(g1762C));
AND2_X1 U_g4903C (.ZN(g4903C),.A2(g4243C),.A1(g1849C));
AND2_X1 U_g11178C (.ZN(g11178C),.A2(FE_OFN13_g10702C),.A1(g516C));
AND2_X1 U_g8510C (.ZN(g8510C),.A2(FE_OFN330_g7638C),.A1(g8414C));
AND2_X1 U_g8245C (.ZN(g8245C),.A2(FE_OFN322_g4449C),.A1(g7062C));
AND2_X1 U_g6319C (.ZN(g6319C),.A2(FE_OFN118_g4807C),.A1(g1296C));
AND2_X1 U_g11186C (.ZN(g11186C),.A2(FE_OFN10_g10702C),.A1(g4722C));
AND2_X1 U_g2951C (.ZN(g2951C),.A2(g1681C),.A1(FE_OFN241_g1690C));
AND2_X1 U_g6352C (.ZN(g6352C),.A2(FE_OFN319_g5361C),.A1(g278C));
AND2_X1 U_g9595C (.ZN(g9595C),.A2(FE_OFN42_g9205C),.A1(g901C));
AND2_X1 U_g4831C (.ZN(g4831C),.A2(g4109C),.A1(g810C));
AND2_X1 U_g5492C (.ZN(g5492C),.A2(g4263C),.A1(g1654C));
AND2_X1 U_g9272C (.ZN(g9272C),.A2(FE_OFN266_g18C),.A1(g8934C));
AND2_X1 U_g10312C (.ZN(g10312C),.A2(g9082C),.A1(g10019C));
AND2_X1 U_g6186C (.ZN(g6186C),.A2(FE_OFN291_g4880C),.A1(g546C));
AND2_X1 U_g9612C (.ZN(g9612C),.A2(FE_OFN40_g9240C),.A1(g2652C));
AND2_X1 U_g9417C (.ZN(g9417C),.A2(FE_OFN56_g9052C),.A1(g1738C));
AND2_X1 U_g9935C (.ZN(g9935C),.A2(FE_OFN60_g9624C),.A1(g9914C));
AND2_X1 U_g10745C (.ZN(g10745C),.A2(FE_OFN102_g3586C),.A1(g10658C));
AND2_X1 U_g11216C (.ZN(g11216C),.A2(FE_OFN279_g11157C),.A1(g956C));
AND2_X1 U_g9328C (.ZN(g9328C),.A2(FE_OFN275_g48C),.A1(g8971C));
AND2_X1 U_g11587C (.ZN(g11587C),.A2(g11539C),.A1(g1327C));
AND2_X1 U_g6821C (.ZN(g6821C),.A2(FE_OFN178_g5354C),.A1(g237C));
AND2_X1 U_g6325C (.ZN(g6325C),.A2(FE_OFN116_g4807C),.A1(g1245C));
AND2_X1 U_g4560C (.ZN(g4560C),.A2(g4002C),.A1(g431C));
AND2_X1 U_g7368C (.ZN(g7368C),.A2(g3880C),.A1(g5842C));
AND2_X1 U_g6083C (.ZN(g6083C),.A2(g4273C),.A1(g552C));
AND2_X1 U_g6544C (.ZN(g6544C),.A2(g6081C),.A1(g1227C));
AND2_X1 U_g5476C (.ZN(g5476C),.A2(g4673C),.A1(g1615C));
AND2_X1 U_g7743C (.ZN(g7743C),.A2(FE_OFN226_g3880C),.A1(g5838C));
AND2_X1 U_g4869C (.ZN(g4869C),.A2(FE_OFN132_g3015C),.A1(g1083C));
AND2_X1 U_g5722C (.ZN(g5722C),.A2(FE_OFN315_g5117C),.A1(g1598C));
AND2_X1 U_g6790C (.ZN(g6790C),.A2(FE_OFN346_g4381C),.A1(g5813C));
AND2_X1 U_g8408C (.ZN(g8408C),.A2(g8146C),.A1(g704C));
AND2_X1 U_g10761C (.ZN(g10761C),.A2(g10558C),.A1(g10559C));
AND2_X1 U_g7734C (.ZN(g7734C),.A2(FE_OFN226_g3880C),.A1(g5810C));
AND2_X1 U_g8136C (.ZN(g8136C),.A2(g7045C),.A1(g7926C));
AND2_X1 U_g6187C (.ZN(g6187C),.A2(g2340C),.A1(g5569C));
AND2_X1 U_g4752C (.ZN(g4752C),.A2(FE_OFN300_g4002C),.A1(g401C));
AND2_X1 U_g9902C (.ZN(g9902C),.A2(FE_OFN69_g9392C),.A1(g9720C));
AND2_X1 U_g8768C (.ZN(g8768C),.A2(FE_OFN304_g5151C),.A1(g8623C));
AND2_X1 U_g5500C (.ZN(g5500C),.A2(g4281C),.A1(g1657C));
AND2_X1 U_g2496C (.ZN(g2496C),.A2(g369C),.A1(g374C));
AND2_X1 U_g6756C (.ZN(g6756C),.A2(g5877C),.A1(g3010C));
AND3_X1 U_g8972C (.ZN(g8972C),.A3(FE_OFN73_g8858C),.A2(FE_OFN281_g2216C),.A1(g8085C));
AND2_X1 U_g6622C (.ZN(g6622C),.A2(g6165C),.A1(g336C));
AND2_X1 U_g11639C (.ZN(g11639C),.A2(g7897C),.A1(g11612C));
AND2_X1 U_g9366C (.ZN(g9366C),.A2(FE_OFN53_g9173C),.A1(g1311C));
AND2_X1 U_g11230C (.ZN(g11230C),.A2(g11060C),.A1(g471C));
AND2_X1 U_g10328C (.ZN(g10328C),.A2(FE_OFN269_g109C),.A1(I15507C));
AND2_X1 U_g5024C (.ZN(g5024C),.A2(FE_OFN303_g4678C),.A1(g1284C));
AND2_X1 U_g4364C (.ZN(g4364C),.A2(g4679C),.A1(g1215C));
AND2_X1 U_g9649C (.ZN(g9649C),.A2(g9205C),.A1(g916C));
AND2_X1 U_g5795C (.ZN(g5795C),.A2(g5261C),.A1(g1543C));
AND2_X1 U_g5737C (.ZN(g5737C),.A2(FE_OFN321_g5261C),.A1(g1524C));
AND2_X1 U_g6841C (.ZN(g6841C),.A2(FE_OFN180_g5354C),.A1(g1400C));
AND2_X1 U_g4054C (.ZN(g4054C),.A2(g2774C),.A1(g1753C));
AND2_X1 U_g6345C (.ZN(g6345C),.A2(FE_OFN346_g4381C),.A1(g5823C));
AND2_X1 U_g11391C (.ZN(g11391C),.A2(g7914C),.A1(g11275C));
AND2_X1 U_g9851C (.ZN(g9851C),.A2(g9764C),.A1(g296C));
AND2_X1 U_g6763C (.ZN(g6763C),.A2(g4381C),.A1(g5802C));
AND2_X1 U_g4770C (.ZN(g4770C),.A2(FE_OFN300_g4002C),.A1(g416C));
AND3_X1 U_I16142C (.ZN(I16142C),.A3(g10507C),.A2(g10509C),.A1(g10511C));
AND2_X1 U_g9698C (.ZN(g9698C),.A2(FE_OFN63_g9474C),.A1(g1571C));
AND2_X1 U_g4725C (.ZN(g4725C),.A2(FE_OFN347_g3914C),.A1(g1032C));
AND2_X1 U_g5477C (.ZN(g5477C),.A2(FE_OFN333_g4294C),.A1(g1887C));
AND2_X1 U_g9964C (.ZN(g9964C),.A2(g9536C),.A1(g9954C));
AND2_X1 U_g5523C (.ZN(g5523C),.A2(g4290C),.A1(g1663C));
AND2_X1 U_g4553C (.ZN(g4553C),.A2(g4002C),.A1(g435C));
AND2_X1 U_g8550C (.ZN(g8550C),.A2(FE_OFN330_g7638C),.A1(g8402C));
AND2_X1 U_g8845C (.ZN(g8845C),.A2(FE_OFN328_g8709C),.A1(g8611C));
AND2_X1 U_g2081C (.ZN(g2081C),.A2(g928C),.A1(g932C));
AND2_X1 U_g6359C (.ZN(g6359C),.A2(FE_OFN320_g5361C),.A1(g281C));
AND2_X1 U_g11586C (.ZN(g11586C),.A2(g11539C),.A1(g1324C));
AND2_X1 U_g11007C (.ZN(g11007C),.A2(FE_OFN13_g10702C),.A1(g5147C));
AND2_X1 U_g5104C (.ZN(g5104C),.A2(g4608C),.A1(g1796C));
AND2_X1 U_g5099C (.ZN(g5099C),.A2(FE_OFN141_g3829C),.A1(g4821C));
AND2_X1 U_g6757C (.ZN(g6757C),.A2(g5919C),.A1(g143C));
AND2_X1 U_g5499C (.ZN(g5499C),.A2(g4679C),.A1(g1627C));
AND2_X1 U_g4389C (.ZN(g4389C),.A2(g3092C),.A1(g3529C));
AND2_X1 U_g6416C (.ZN(g6416C),.A2(FE_OFN217_g5013C),.A1(g3497C));
AND2_X1 U_g9720C (.ZN(g9720C),.A2(g9490C),.A1(g1546C));
AND2_X1 U_g4990C (.ZN(g4990C),.A2(FE_OFN147_g4682C),.A1(g1444C));
AND2_X1 U_g9619C (.ZN(g9619C),.A2(g9010C),.A1(g940C));
AND4_X1 U_I6630C (.ZN(I6630C),.A4(FE_OFN253_g1786C),.A3(FE_OFN236_g1776C),.A2(FE_OFN247_g1771C),.A1(g2677C));
AND2_X1 U_g6047C (.ZN(g6047C),.A2(g4977C),.A1(g2017C));
AND2_X1 U_g9652C (.ZN(g9652C),.A2(FE_OFN39_g9223C),.A1(g953C));
AND3_X1 U_g10515C (.ZN(g10515C),.A3(I16142C),.A2(g10469C),.A1(g10505C));
AND2_X1 U_g9843C (.ZN(g9843C),.A2(g9519C),.A1(g9711C));
AND2_X1 U_g5273C (.ZN(g5273C),.A2(g4776C),.A1(g1074C));
AND2_X1 U_g11465C (.ZN(g11465C),.A2(FE_OFN100_g4421C),.A1(g11232C));
AND2_X1 U_g5044C (.ZN(g5044C),.A2(g1918C),.A1(g4348C));
AND2_X1 U_g11237C (.ZN(g11237C),.A2(g11111C),.A1(g4548C));
AND2_X1 U_g9834C (.ZN(g9834C),.A2(FE_OFN34_g9785C),.A1(g9731C));
AND2_X1 U_g6654C (.ZN(g6654C),.A2(FE_OFN282_g6165C),.A1(g363C));
AND2_X1 U_g5444C (.ZN(g5444C),.A2(FE_OFN290_g4880C),.A1(g1041C));
AND2_X1 U_g3714C (.ZN(g3714C),.A2(g2299C),.A1(g1690C));
AND2_X1 U_g11340C (.ZN(g11340C),.A2(g4285C),.A1(g11285C));
AND2_X1 U_g9598C (.ZN(g9598C),.A2(g9274C),.A1(g119C));
AND2_X1 U_g8097C (.ZN(g8097C),.A2(g7852C),.A1(g5477C));
AND2_X1 U_g8726C (.ZN(g8726C),.A2(g7913C),.A1(g8221C));
AND2_X1 U_g6880C (.ZN(g6880C),.A2(g6557C),.A1(g4816C));
AND2_X1 U_g4338C (.ZN(g4338C),.A2(FE_OFN351_g3913C),.A1(g1157C));
AND2_X1 U_g5543C (.ZN(g5543C),.A2(FE_OFN322_g4449C),.A1(g2979C));
AND3_X1 U_g8960C (.ZN(g8960C),.A3(g8828C),.A2(FE_OFN95_g2216C),.A1(g8085C));
AND2_X1 U_g4109C (.ZN(g4109C),.A2(g3287C),.A1(g806C));
AND2_X1 U_g10759C (.ZN(g10759C),.A2(g10556C),.A1(g10557C));
AND2_X1 U_g9938C (.ZN(g9938C),.A2(FE_OFN67_g9367C),.A1(g9917C));
AND2_X1 U_g10758C (.ZN(g10758C),.A2(FE_OFN293_g3015C),.A1(g10652C));
AND2_X1 U_g4759C (.ZN(g4759C),.A2(FE_OFN300_g4002C),.A1(g406C));
AND2_X1 U_g9909C (.ZN(g9909C),.A2(FE_OFN33_g9454C),.A1(g9891C));
AND2_X1 U_g7127C (.ZN(g7127C),.A2(g2241C),.A1(g6663C));
AND2_X1 U_g11165C (.ZN(g11165C),.A2(FE_OFN13_g10702C),.A1(g476C));
AND2_X1 U_g6234C (.ZN(g6234C),.A2(FE_OFN306_g5128C),.A1(g1424C));
AND2_X1 U_g6328C (.ZN(g6328C),.A2(FE_OFN115_g4807C),.A1(g1260C));
AND2_X1 U_g8401C (.ZN(g8401C),.A2(g8146C),.A1(g677C));
AND2_X1 U_g11006C (.ZN(g11006C),.A2(FE_OFN18_g10702C),.A1(g5125C));
AND2_X1 U_g4865C (.ZN(g4865C),.A2(FE_OFN297_g3015C),.A1(g1080C));
AND2_X1 U_g4715C (.ZN(g4715C),.A2(FE_OFN297_g3015C),.A1(g1077C));
AND3_X1 U_g4604C (.ZN(g4604C),.A3(g2325C),.A2(g3753C),.A1(g3056C));
AND2_X1 U_g5513C (.ZN(g5513C),.A2(g3906C),.A1(g1675C));
AND2_X1 U_g11222C (.ZN(g11222C),.A2(FE_OFN279_g11157C),.A1(g965C));
AND2_X1 U_g4498C (.ZN(g4498C),.A2(FE_OFN302_g3913C),.A1(g1145C));
AND2_X1 U_g6554C (.ZN(g6554C),.A2(g5808C),.A1(g96C));
AND2_X1 U_g7732C (.ZN(g7732C),.A2(FE_OFN226_g3880C),.A1(g5803C));
AND2_X1 U_g9586C (.ZN(g9586C),.A2(FE_OFN53_g9173C),.A1(g1346C));
AND3_X1 U_g5178C (.ZN(g5178C),.A3(g4104C),.A2(FE_OFN223_g4401C),.A1(g2047C));
AND2_X1 U_g4584C (.ZN(g4584C),.A2(g1857C),.A1(g3710C));
AND2_X1 U_g7472C (.ZN(g7472C),.A2(g61C),.A1(FE_OFN83_g2176C));
AND2_X1 U_g11253C (.ZN(g11253C),.A2(g11083C),.A1(g981C));
AND2_X1 U_g5182C (.ZN(g5182C),.A2(FE_OFN303_g4678C),.A1(g1240C));
AND2_X1 U_g9860C (.ZN(g9860C),.A2(g9778C),.A1(g1598C));
AND2_X1 U_g11600C (.ZN(g11600C),.A2(g11575C),.A1(g1346C));
AND2_X1 U_g9710C (.ZN(g9710C),.A2(FE_OFN63_g9474C),.A1(g1586C));
AND2_X1 U_g9645C (.ZN(g9645C),.A2(FE_OFN51_g9111C),.A1(g1203C));
AND2_X1 U_g11236C (.ZN(g11236C),.A2(g11111C),.A1(g4537C));
AND2_X1 U_g4162C (.ZN(g4162C),.A2(g1845C),.A1(g3106C));
AND2_X1 U_g6090C (.ZN(g6090C),.A2(g5627C),.A1(g553C));
AND2_X1 U_g9691C (.ZN(g9691C),.A2(g9432C),.A1(g269C));
AND2_X1 U_g11372C (.ZN(g11372C),.A2(g4285C),.A1(g11316C));
AND2_X1 U_g6823C (.ZN(g6823C),.A2(g5354C),.A1(g1368C));
AND2_X1 U_g11175C (.ZN(g11175C),.A2(FE_OFN20_g10702C),.A1(g501C));
AND2_X1 U_g8068C (.ZN(g8068C),.A2(FE_OFN198_g7697C),.A1(g664C));
AND2_X1 U_g9607C (.ZN(g9607C),.A2(g9274C),.A1(g12C));
AND2_X1 U_g9962C (.ZN(g9962C),.A2(FE_OFN280_g9536C),.A1(g9952C));
AND2_X1 U_g6348C (.ZN(g6348C),.A2(FE_OFN320_g5361C),.A1(g296C));
AND2_X1 U_g9659C (.ZN(g9659C),.A2(FE_OFN39_g9223C),.A1(g956C));
AND2_X1 U_g9358C (.ZN(g9358C),.A2(FE_OFN47_g9151C),.A1(g1318C));
AND2_X1 U_g3104C (.ZN(g3104C),.A2(I6317C),.A1(I6316C));
AND2_X1 U_g4486C (.ZN(g4486C),.A2(g4679C),.A1(g1711C));
AND2_X1 U_g9587C (.ZN(g9587C),.A2(g8995C),.A1(g892C));
AND2_X1 U_g5632C (.ZN(g5632C),.A2(I5435C),.A1(g1636C));
AND2_X4 U_g9111C (.ZN(g9111C),.A2(FE_OFN276_g48C),.A1(g8965C));
AND2_X1 U_g4881C (.ZN(g4881C),.A2(FE_OFN347_g3914C),.A1(g991C));
AND2_X1 U_g11209C (.ZN(g11209C),.A2(FE_OFN79_g8700C),.A1(g10712C));
AND2_X1 U_g8848C (.ZN(g8848C),.A2(FE_OFN328_g8709C),.A1(g8715C));
AND2_X1 U_g4070C (.ZN(g4070C),.A2(g2330C),.A1(g3263C));
AND2_X1 U_g6463C (.ZN(g6463C),.A2(I9237C),.A1(FE_OFN277_g48C));
AND4_X1 U_I5689C (.ZN(I5689C),.A4(g1432C),.A3(g1428C),.A2(g1424C),.A1(g1419C));
AND2_X1 U_g7820C (.ZN(g7820C),.A2(FE_OFN209_g6863C),.A1(g1896C));
AND2_X1 U_g11021C (.ZN(g11021C),.A2(FE_OFN7_g10702C),.A1(g448C));
AND2_X1 U_g5917C (.ZN(g5917C),.A2(g85C),.A1(g1044C));
AND2_X1 U_g6619C (.ZN(g6619C),.A2(FE_OFN97_I8869C),.A1(g49C));
AND2_X1 U_g6318C (.ZN(g6318C),.A2(FE_OFN118_g4807C),.A1(g1300C));
AND2_X1 U_g6872C (.ZN(g6872C),.A2(FE_OFN213_g6003C),.A1(g1896C));
AND2_X1 U_g11320C (.ZN(g11320C),.A2(g4379C),.A1(g11201C));
AND2_X1 U_g10514C (.ZN(g10514C),.A2(FE_OFN370_g4525C),.A1(g10489C));
AND2_X1 U_g4006C (.ZN(g4006C),.A2(FE_OFN266_g18C),.A1(g201C));
AND2_X1 U_g9853C (.ZN(g9853C),.A2(g9764C),.A1(g299C));
AND2_X1 U_g11274C (.ZN(g11274C),.A2(g11199C),.A1(g4771C));
AND2_X1 U_g6193C (.ZN(g6193C),.A2(FE_OFN306_g5128C),.A1(g1419C));
AND2_X1 U_g8119C (.ZN(g8119C),.A2(FE_OFN207_g6863C),.A1(g5526C));
AND2_X1 U_g9420C (.ZN(g9420C),.A2(FE_OFN50_g9030C),.A1(g1747C));
AND2_X1 U_g5233C (.ZN(g5233C),.A2(g4492C),.A1(FE_OFN252_g1791C));
AND2_X1 U_g7581C (.ZN(g7581C),.A2(g5420C),.A1(g7092C));
AND2_X1 U_g6549C (.ZN(g6549C),.A2(g5808C),.A1(g95C));
AND2_X1 U_g11464C (.ZN(g11464C),.A2(FE_OFN100_g4421C),.A1(g11231C));
AND2_X1 U_g4801C (.ZN(g4801C),.A2(FE_OFN307_g4010C),.A1(g516C));
AND2_X1 U_g6834C (.ZN(g6834C),.A2(FE_OFN178_g5354C),.A1(g1365C));
AND2_X1 U_g4487C (.ZN(g4487C),.A2(g3906C),.A1(g1718C));
AND2_X1 U_g2939C (.ZN(g2939C),.A2(g1687C),.A1(FE_OFN241_g1690C));
AND2_X1 U_g7060C (.ZN(g7060C),.A2(g5521C),.A1(g6739C));
AND2_X1 U_g5770C (.ZN(g5770C),.A2(g5128C),.A1(g3585C));
AND2_X1 U_g5725C (.ZN(g5725C),.A2(FE_OFN353_g5117C),.A1(g1580C));
AND2_X1 U_g11641C (.ZN(g11641C),.A2(g7897C),.A1(g11615C));
AND2_X1 U_g2544C (.ZN(g2544C),.A2(g1336C),.A1(g1341C));
AND2_X1 U_g11292C (.ZN(g11292C),.A2(g4379C),.A1(g11252C));
AND2_X1 U_g5532C (.ZN(g5532C),.A2(g4273C),.A1(g1681C));
AND2_X1 U_g11153C (.ZN(g11153C),.A2(g10788C),.A1(g3771C));
AND2_X1 U_g9905C (.ZN(g9905C),.A2(g9680C),.A1(g9872C));
AND2_X1 U_g7739C (.ZN(g7739C),.A2(g3880C),.A1(g5820C));
AND2_X1 U_g6321C (.ZN(g6321C),.A2(FE_OFN118_g4807C),.A1(g1284C));
AND2_X1 U_g8386C (.ZN(g8386C),.A2(g8220C),.A1(g5257C));
AND3_X1 U_g8975C (.ZN(g8975C),.A3(FE_OFN73_g8858C),.A2(FE_OFN281_g2216C),.A1(g8089C));
AND2_X1 U_g2306C (.ZN(g2306C),.A2(g1218C),.A1(g1223C));
AND2_X1 U_g6625C (.ZN(g6625C),.A2(g6081C),.A1(g1218C));
AND2_X1 U_g7937C (.ZN(g7937C),.A2(FE_OFN292_g3015C),.A1(g5274C));
AND2_X2 U_g10788C (.ZN(g10788C),.A2(g10702C),.A1(g8303C));
AND2_X1 U_g10325C (.ZN(g10325C),.A2(FE_OFN352_g109C),.A1(I15503C));
AND2_X1 U_g8170C (.ZN(g8170C),.A2(FE_OFN89_I11360C),.A1(g36C));
AND2_X1 U_g5706C (.ZN(g5706C),.A2(FE_OFN315_g5117C),.A1(g1574C));
AND2_X1 U_g2756C (.ZN(g2756C),.A2(g2081C),.A1(g936C));
AND2_X1 U_g8821C (.ZN(g8821C),.A2(FE_OFN328_g8709C),.A1(g8643C));
AND2_X1 U_g10946C (.ZN(g10946C),.A2(FE_OFN9_g10702C),.A1(g5225C));
AND2_X1 U_g4169C (.ZN(g4169C),.A2(g3060C),.A1(FE_OFN237_g1806C));
AND2_X1 U_g5029C (.ZN(g5029C),.A2(FE_OFN288_g4263C),.A1(g1077C));
AND2_X1 U_g11164C (.ZN(g11164C),.A2(FE_OFN13_g10702C),.A1(g3513C));
AND2_X1 U_g4007C (.ZN(g4007C),.A2(g2276C),.A1(FE_OFN247_g1771C));
AND2_X1 U_g4059C (.ZN(g4059C),.A2(g2774C),.A1(g1756C));
AND2_X1 U_g4868C (.ZN(g4868C),.A2(FE_OFN347_g3914C),.A1(g1027C));
AND2_X1 U_g5675C (.ZN(g5675C),.A2(FE_OFN365_g5361C),.A1(g131C));
AND2_X1 U_g4718C (.ZN(g4718C),.A2(g3943C),.A1(g650C));
AND2_X1 U_g10682C (.ZN(g10682C),.A2(FE_OFN136_g3863C),.A1(g10381C));
AND2_X1 U_g6687C (.ZN(g6687C),.A2(I9326C),.A1(g92C));
AND2_X1 U_g7704C (.ZN(g7704C),.A2(FE_OFN191_g6488C),.A1(g682C));
AND2_X1 U_g4582C (.ZN(g4582C),.A2(g4010C),.A1(g525C));
AND2_X1 U_g4261C (.ZN(g4261C),.A2(FE_OFN347_g3914C),.A1(g1019C));
AND2_X1 U_g3422C (.ZN(g3422C),.A2(FE_OFN324_g18C),.A1(g225C));
AND2_X1 U_g5745C (.ZN(g5745C),.A2(FE_OFN321_g5261C),.A1(g1549C));
AND2_X1 U_g8387C (.ZN(g8387C),.A2(g8220C),.A1(g5258C));
AND2_X1 U_g7954C (.ZN(g7954C),.A2(g7512C),.A1(g49C));
AND2_X1 U_g11283C (.ZN(g11283C),.A2(g11239C),.A1(g4804C));
AND2_X1 U_g8461C (.ZN(g8461C),.A2(FE_OFN210_g7246C),.A1(g8298C));
AND2_X1 U_g10760C (.ZN(g10760C),.A2(g10554C),.A1(g10555C));
AND2_X1 U_g11492C (.ZN(g11492C),.A2(g4807C),.A1(g11480C));
AND3_X1 U_g7032C (.ZN(g7032C),.A3(I7048C),.A2(g6626C),.A1(g109C));
AND2_X4 U_g9151C (.ZN(g9151C),.A2(FE_OFN276_g48C),.A1(g8967C));
AND2_X1 U_g6341C (.ZN(g6341C),.A2(FE_OFN319_g5361C),.A1(g272C));
AND2_X1 U_g10506C (.ZN(g10506C),.A2(FE_OFN241_g1690C),.A1(g10007C));
AND2_X1 U_g9648C (.ZN(g9648C),.A2(FE_OFN62_g9274C),.A1(g16C));
AND2_X1 U_g7453C (.ZN(g7453C),.A2(g52C),.A1(FE_OFN86_g2176C));
AND2_X1 U_g6525C (.ZN(g6525C),.A2(FE_OFN343_I5565C),.A1(g5995C));
AND2_X1 U_g6645C (.ZN(g6645C),.A2(FE_OFN97_I8869C),.A1(g67C));
AND2_X1 U_g5707C (.ZN(g5707C),.A2(FE_OFN353_g5117C),.A1(g1595C));
AND2_X1 U_g8046C (.ZN(g8046C),.A2(FE_OFN305_g5151C),.A1(g7548C));
AND2_X1 U_g11091C (.ZN(g11091C),.A2(FE_OFN4_g10950C),.A1(g833C));
AND2_X1 U_g11174C (.ZN(g11174C),.A2(FE_OFN21_g10702C),.A1(g496C));
AND2_X4 U_g9010C (.ZN(g9010C),.A2(g8930C),.A1(FE_OFN277_g48C));
AND2_X1 U_g8403C (.ZN(g8403C),.A2(g8220C),.A1(g5276C));
AND2_X1 U_g5201C (.ZN(g5201C),.A2(g4678C),.A1(g1250C));
AND2_X1 U_g8841C (.ZN(g8841C),.A2(FE_OFN328_g8709C),.A1(g8605C));
AND2_X1 U_g6879C (.ZN(g6879C),.A2(FE_OFN213_g6003C),.A1(g1914C));
AND2_X2 U_g8763C (.ZN(g8763C),.A2(g8451C),.A1(I9880C));
AND2_X1 U_g4502C (.ZN(g4502C),.A2(g3938C),.A1(g2031C));
AND2_X1 U_g9839C (.ZN(g9839C),.A2(g9747C),.A1(g9702C));
AND2_X1 U_g6358C (.ZN(g6358C),.A2(FE_OFN346_g4381C),.A1(g5841C));
AND2_X1 U_g5575C (.ZN(g5575C),.A2(FE_OFN367_g3521C),.A1(g1618C));
AND2_X1 U_g4940C (.ZN(g4940C),.A2(FE_OFN310_g4336C),.A1(g1984C));
AND2_X1 U_g8107C (.ZN(g8107C),.A2(g7852C),.A1(g5502C));
AND2_X1 U_g10240C (.ZN(g10240C),.A2(g9082C),.A1(g9974C));
AND2_X1 U_g11192C (.ZN(g11192C),.A2(g10927C),.A1(g4759C));
AND2_X1 U_g9618C (.ZN(g9618C),.A2(g9205C),.A1(g910C));
AND2_X1 U_g5539C (.ZN(g5539C),.A2(g4273C),.A1(g1684C));
AND2_X1 U_g8416C (.ZN(g8416C),.A2(FE_OFN187_g7638C),.A1(g731C));
AND2_X1 U_g9693C (.ZN(g9693C),.A2(FE_OFN59_g9432C),.A1(g275C));
AND2_X1 U_g11553C (.ZN(g11553C),.A2(g11519C),.A1(g1771C));
AND2_X1 U_g8047C (.ZN(g8047C),.A2(FE_OFN177_g5919C),.A1(g7557C));
AND2_X1 U_g5268C (.ZN(g5268C),.A2(g4263C),.A1(g1098C));
AND2_X1 U_g9555C (.ZN(g9555C),.A2(FE_OFN325_g18C),.A1(g9107C));
AND2_X1 U_g6180C (.ZN(g6180C),.A2(g5128C),.A1(g1453C));
AND2_X1 U_g6832C (.ZN(g6832C),.A2(FE_OFN179_g5354C),.A1(g1383C));
AND2_X1 U_g10633C (.ZN(g10633C),.A2(g3829C),.A1(g10381C));
AND2_X1 U_g7894C (.ZN(g7894C),.A2(FE_OFN366_g3521C),.A1(g5317C));
AND2_X1 U_g8654C (.ZN(g8654C),.A2(FE_OFN348_g3015C),.A1(g8266C));
AND2_X1 U_g9621C (.ZN(g9621C),.A2(FE_OFN46_g9125C),.A1(g1179C));
AND2_X1 U_g6794C (.ZN(g6794C),.A2(FE_OFN346_g4381C),.A1(g5819C));
AND2_X1 U_g9313C (.ZN(g9313C),.A2(FE_OFN275_g48C),.A1(g8876C));
AND2_X1 U_g3412C (.ZN(g3412C),.A2(g18C),.A1(g219C));
AND2_X1 U_g7661C (.ZN(g7661C),.A2(g2251C),.A1(g7127C));
AND3_X1 U_g2800C (.ZN(g2800C),.A3(g591C),.A2(g2369C),.A1(g2399C));
AND2_X1 U_g3706C (.ZN(g3706C),.A2(g3268C),.A1(g471C));
AND2_X1 U_g9908C (.ZN(g9908C),.A2(FE_OFN33_g9454C),.A1(g9760C));
AND2_X1 U_g3429C (.ZN(g3429C),.A2(g18C),.A1(g231C));
AND2_X1 U_g6628C (.ZN(g6628C),.A2(FE_OFN282_g6165C),.A1(g351C));
AND2_X1 U_g5470C (.ZN(g5470C),.A2(g4880C),.A1(g1044C));
AND2_X1 U_g7526C (.ZN(g7526C),.A2(g73C),.A1(FE_OFN87_g2176C));
AND2_X1 U_g5897C (.ZN(g5897C),.A2(g5354C),.A1(g2204C));
AND2_X1 U_g5025C (.ZN(g5025C),.A2(FE_OFN153_g4640C),.A1(g1482C));
AND2_X1 U_g6204C (.ZN(g6204C),.A2(FE_OFN200_g4921C),.A1(g3738C));
AND2_X1 U_g4048C (.ZN(g4048C),.A2(g2774C),.A1(g1750C));
AND3_X1 U_g8935C (.ZN(g8935C),.A3(g8849C),.A2(FE_OFN95_g2216C),.A1(g8106C));
AND2_X1 U_g3281C (.ZN(g3281C),.A2(g2525C),.A1(g766C));
AND2_X1 U_g9593C (.ZN(g9593C),.A2(FE_OFN42_g9205C),.A1(g898C));
AND2_X1 U_g4827C (.ZN(g4827C),.A2(FE_OFN324_g18C),.A1(g213C));
AND2_X1 U_g10701C (.ZN(g10701C),.A2(g10500C),.A1(g10501C));
AND2_X1 U_g10777C (.ZN(g10777C),.A2(g3015C),.A1(g10733C));
AND2_X1 U_g8130C (.ZN(g8130C),.A2(g7952C),.A1(g1936C));
AND2_X1 U_g9965C (.ZN(g9965C),.A2(FE_OFN280_g9536C),.A1(g9955C));
AND2_X1 U_g3684C (.ZN(g3684C),.A2(g3015C),.A1(g1710C));
AND2_X1 U_g11213C (.ZN(g11213C),.A2(FE_OFN279_g11157C),.A1(g947C));
AND2_X1 U_g5006C (.ZN(g5006C),.A2(FE_OFN154_g4640C),.A1(g1462C));
AND2_X1 U_g9933C (.ZN(g9933C),.A2(g9624C),.A1(g9912C));
AND2_X1 U_g8554C (.ZN(g8554C),.A2(FE_OFN330_g7638C),.A1(g8407C));
AND2_X1 U_g9641C (.ZN(g9641C),.A2(g9205C),.A1(g913C));
AND2_X1 U_g6123C (.ZN(g6123C),.A2(FE_OFN310_g4336C),.A1(g3662C));
AND2_X1 U_g6323C (.ZN(g6323C),.A2(FE_OFN116_g4807C),.A1(g1235C));
AND2_X1 U_g10766C (.ZN(g10766C),.A2(FE_OFN131_g3015C),.A1(g10646C));
AND2_X1 U_g6666C (.ZN(g6666C),.A2(g5836C),.A1(g89C));
AND2_X1 U_g4994C (.ZN(g4994C),.A2(FE_OFN154_g4640C),.A1(g1504C));
AND2_X1 U_g5755C (.ZN(g5755C),.A2(FE_OFN179_g5354C),.A1(g5103C));
AND2_X1 U_g11592C (.ZN(g11592C),.A2(g11561C),.A1(g3717C));
AND2_X1 U_g6351C (.ZN(g6351C),.A2(g48C),.A1(I9237C));
AND2_X1 U_g6875C (.ZN(g6875C),.A2(FE_OFN213_g6003C),.A1(g1905C));
AND2_X1 U_g4816C (.ZN(g4816C),.A2(g2336C),.A1(g4070C));
AND2_X1 U_g9658C (.ZN(g9658C),.A2(g9240C),.A1(g947C));
AND2_X1 U_g6530C (.ZN(g6530C),.A2(FE_OFN141_g3829C),.A1(g6207C));
AND2_X1 U_g8366C (.ZN(g8366C),.A2(g7265C),.A1(g8199C));
AND2_X1 U_g9835C (.ZN(g9835C),.A2(FE_OFN34_g9785C),.A1(g9735C));
AND2_X1 U_g6655C (.ZN(g6655C),.A2(I9326C),.A1(g88C));
AND3_X1 U_g5445C (.ZN(g5445C),.A3(g109C),.A2(g3875C),.A1(FE_OFN184_I7048C));
AND2_X1 U_g5173C (.ZN(g5173C),.A2(g4671C),.A1(g1110C));
AND2_X1 U_g7970C (.ZN(g7970C),.A2(g7438C),.A1(g7384C));
AND2_X1 U_g3098C (.ZN(g3098C),.A2(g2198C),.A1(g2331C));
AND2_X1 U_g5491C (.ZN(g5491C),.A2(g4289C),.A1(g1624C));
AND2_X1 U_g9271C (.ZN(g9271C),.A2(g8949C),.A1(g6109C));
AND2_X1 U_g11152C (.ZN(g11152C),.A2(g10883C),.A1(g369C));
AND2_X1 U_g9611C (.ZN(g9611C),.A2(g9010C),.A1(g936C));
AND2_X1 U_g6410C (.ZN(g6410C),.A2(FE_OFN217_g5013C),.A1(g2804C));
AND2_X1 U_g10451C (.ZN(g10451C),.A2(g2024C),.A1(g10444C));
AND2_X1 U_g4397C (.ZN(g4397C),.A2(g639C),.A1(g3475C));
AND2_X1 U_g7224C (.ZN(g7224C),.A2(g6447C),.A1(g5398C));
AND2_X1 U_g5602C (.ZN(g5602C),.A2(FE_OFN357_g3521C),.A1(g1624C));
AND2_X2 U_g4421C (.ZN(g4421C),.A2(g750C),.A1(g2057C));
AND2_X1 U_g6884C (.ZN(g6884C),.A2(g6557C),.A1(g5569C));
AND2_X1 U_g6839C (.ZN(g6839C),.A2(FE_OFN180_g5354C),.A1(g1397C));
AND3_X1 U_g8964C (.ZN(g8964C),.A3(g8849C),.A2(FE_OFN92_g2216C),.A1(g8255C));
AND2_X1 U_g8260C (.ZN(g8260C),.A2(g7907C),.A1(g940C));
AND2_X1 U_g11413C (.ZN(g11413C),.A2(g10679C),.A1(g11217C));
AND2_X1 U_g4950C (.ZN(g4950C),.A2(FE_OFN146_g4682C),.A1(g1415C));
AND2_X1 U_g5535C (.ZN(g5535C),.A2(FE_OFN366_g3521C),.A1(g572C));
AND2_X1 U_g7277C (.ZN(g7277C),.A2(g731C),.A1(g6772C));
AND2_X1 U_g8463C (.ZN(g8463C),.A2(FE_OFN211_g7246C),.A1(g8301C));
AND2_X1 U_g3268C (.ZN(g3268C),.A2(g2511C),.A1(FE_OFN248_g466C));
AND2_X1 U_g10785C (.ZN(g10785C),.A2(g4467C),.A1(g10728C));
AND2_X1 U_g6618C (.ZN(g6618C),.A2(FE_OFN219_g5557C),.A1(g658C));
AND2_X1 U_g6235C (.ZN(g6235C),.A2(g5613C),.A1(g569C));
AND2_X1 U_g10950C (.ZN(g10950C),.A2(g6355C),.A1(g10788C));
AND2_X1 U_g4723C (.ZN(g4723C),.A2(g627C),.A1(g3626C));
AND2_X1 U_g8720C (.ZN(g8720C),.A2(g7905C),.A1(g8206C));
AND2_X1 U_g6693C (.ZN(g6693C),.A2(I9326C),.A1(g93C));
AND2_X1 U_g11020C (.ZN(g11020C),.A2(FE_OFN7_g10702C),.A1(g452C));
AND2_X1 U_g11583C (.ZN(g11583C),.A2(g11539C),.A1(g1314C));
AND2_X1 U_g8118C (.ZN(g8118C),.A2(g7949C),.A1(g1900C));
AND2_X1 U_g8167C (.ZN(g8167C),.A2(FE_OFN89_I11360C),.A1(g33C));
AND2_X1 U_g6334C (.ZN(g6334C),.A2(FE_OFN180_g5354C),.A1(g1389C));
AND2_X1 U_g7892C (.ZN(g7892C),.A2(g3814C),.A1(g5308C));
AND2_X1 U_g8652C (.ZN(g8652C),.A2(FE_OFN119_g3015C),.A1(g8264C));
AND2_X1 U_g5721C (.ZN(g5721C),.A2(FE_OFN353_g5117C),.A1(g1577C));
AND2_X1 U_g10367C (.ZN(g10367C),.A2(FE_OFN234_g2024C),.A1(g10362C));
AND2_X1 U_g9901C (.ZN(g9901C),.A2(FE_OFN69_g9392C),.A1(g9719C));
AND2_X1 U_g6792C (.ZN(g6792C),.A2(FE_OFN319_g5361C),.A1(g290C));
AND2_X1 U_g11282C (.ZN(g11282C),.A2(g11203C),.A1(g4801C));
AND2_X1 U_g7945C (.ZN(g7945C),.A2(g7473C),.A1(g67C));
AND3_X1 U_g8971C (.ZN(g8971C),.A3(FE_OFN73_g8858C),.A2(FE_OFN281_g2216C),.A1(g8081C));
AND2_X1 U_g11302C (.ZN(g11302C),.A2(g11243C),.A1(g4582C));
AND2_X1 U_g4585C (.ZN(g4585C),.A2(g4010C),.A1(g521C));
AND2_X1 U_g6621C (.ZN(g6621C),.A2(I8869C),.A1(g52C));
AND2_X1 U_g5502C (.ZN(g5502C),.A2(FE_OFN333_g4294C),.A1(g1932C));
AND2_X1 U_g11105C (.ZN(g11105C),.A2(g10937C),.A1(g3634C));
AND2_X1 U_g7709C (.ZN(g7709C),.A2(FE_OFN322_g4449C),.A1(g5942C));
AND2_X1 U_g8598C (.ZN(g8598C),.A2(FE_OFN210_g7246C),.A1(g8471C));
AND2_X1 U_g7140C (.ZN(g7140C),.A2(g6716C),.A1(g5221C));
AND2_X1 U_g9600C (.ZN(g9600C),.A2(FE_OFN42_g9205C),.A1(g904C));
AND2_X1 U_g9864C (.ZN(g9864C),.A2(g9778C),.A1(g1604C));
AND2_X1 U_g11640C (.ZN(g11640C),.A2(g7897C),.A1(g11613C));
AND2_X1 U_g5188C (.ZN(g5188C),.A2(g794C),.A1(g798C));
AND2_X1 U_g7435C (.ZN(g7435C),.A2(g6403C),.A1(g7260C));
AND2_X1 U_g7876C (.ZN(g7876C),.A2(FE_OFN366_g3521C),.A1(g5278C));
AND2_X1 U_g5030C (.ZN(g5030C),.A2(FE_OFN303_g4678C),.A1(g1280C));
AND2_X1 U_g4058C (.ZN(g4058C),.A2(FE_OFN224_g2276C),.A1(FE_OFN252_g1791C));
AND2_X1 U_g6776C (.ZN(g6776C),.A2(FE_OFN111_g3914C),.A1(g5809C));
AND2_X1 U_g4890C (.ZN(g4890C),.A2(g4739C),.A1(g630C));
AND2_X1 U_g2525C (.ZN(g2525C),.A2(g758C),.A1(g762C));
AND2_X1 U_g10301C (.ZN(g10301C),.A2(g10025C),.A1(g8700C));
AND2_X1 U_g4505C (.ZN(g4505C),.A2(FE_OFN287_g3586C),.A1(g354C));
AND2_X1 U_g9623C (.ZN(g9623C),.A2(FE_OFN62_g9274C),.A1(g17C));
AND2_X1 U_g10739C (.ZN(g10739C),.A2(g3368C),.A1(g10676C));
AND2_X1 U_g11027C (.ZN(g11027C),.A2(FE_OFN17_g10702C),.A1(g391C));
AND2_X1 U_g10738C (.ZN(g10738C),.A2(FE_OFN131_g3015C),.A1(g10599C));
AND2_X1 U_g8687C (.ZN(g8687C),.A2(FE_OFN189_g7638C),.A1(g8558C));
AND2_X1 U_g6360C (.ZN(g6360C),.A2(FE_OFN319_g5361C),.A1(g302C));
AND2_X1 U_g9871C (.ZN(g9871C),.A2(g9802C),.A1(g1564C));
AND2_X1 U_g5108C (.ZN(g5108C),.A2(g4608C),.A1(g1801C));
AND2_X1 U_g11248C (.ZN(g11248C),.A2(g11083C),.A1(g976C));
AND2_X1 U_g4992C (.ZN(g4992C),.A2(FE_OFN147_g4682C),.A1(g1407C));
AND2_X1 U_g11552C (.ZN(g11552C),.A2(FE_OFN27_g11519C),.A1(g2677C));
AND2_X1 U_g9651C (.ZN(g9651C),.A2(g9240C),.A1(g944C));
AND2_X1 U_g11204C (.ZN(g11204C),.A2(g11083C),.A1(g971C));
AND2_X1 U_g7824C (.ZN(g7824C),.A2(FE_OFN206_g6863C),.A1(g1932C));
AND2_X1 U_g4480C (.ZN(g4480C),.A2(FE_OFN302_g3913C),.A1(g1133C));
AND2_X1 U_g6179C (.ZN(g6179C),.A2(g5354C),.A1(g5115C));
AND2_X1 U_g7590C (.ZN(g7590C),.A2(g5420C),.A1(g7102C));
AND2_X1 U_g9384C (.ZN(g9384C),.A2(g9223C),.A1(g968C));
AND2_X1 U_g3407C (.ZN(g3407C),.A2(FE_OFN352_g109C),.A1(g2561C));
AND2_X1 U_g9838C (.ZN(g9838C),.A2(g9754C),.A1(g9700C));
AND2_X1 U_g10661C (.ZN(g10661C),.A2(FE_OFN119_g3015C),.A1(g10594C));
AND2_X1 U_g11380C (.ZN(g11380C),.A2(g4285C),.A1(g11321C));
AND3_X1 U_g8879C (.ZN(g8879C),.A3(FE_OFN73_g8858C),.A2(FE_OFN281_g2216C),.A1(g8110C));
AND2_X1 U_g7930C (.ZN(g7930C),.A2(FE_OFN343_I5565C),.A1(g7621C));
AND3_X1 U_g8962C (.ZN(g8962C),.A3(g8828C),.A2(FE_OFN95_g2216C),.A1(g8089C));
AND2_X1 U_g10715C (.ZN(g10715C),.A2(g10584C),.A1(g2272C));
AND2_X1 U_g8659C (.ZN(g8659C),.A2(FE_OFN298_g3015C),.A1(g8269C));
AND2_X4 U_g3015C (.ZN(g3015C),.A2(I6260C),.A1(g2028C));
AND2_X1 U_g9643C (.ZN(g9643C),.A2(FE_OFN39_g9223C),.A1(g950C));
AND2_X4 U_g9205C (.ZN(g9205C),.A2(g8957C),.A1(FE_OFN276_g48C));
AND2_X1 U_g5538C (.ZN(g5538C),.A2(FE_OFN288_g4263C),.A1(g1669C));
AND2_X1 U_g4000C (.ZN(g4000C),.A2(g2774C),.A1(g1744C));
AND2_X1 U_g4126C (.ZN(g4126C),.A2(g3060C),.A1(FE_OFN253_g1786C));
AND2_X1 U_g4400C (.ZN(g4400C),.A2(FE_OFN137_g3829C),.A1(g4088C));
AND2_X1 U_g2794C (.ZN(g2794C),.A2(I5887C),.A1(I5886C));
AND2_X1 U_g4760C (.ZN(g4760C),.A2(FE_OFN307_g4010C),.A1(g486C));
AND2_X1 U_g6238C (.ZN(g6238C),.A2(FE_OFN289_g4679C),.A1(g572C));
AND2_X1 U_g10784C (.ZN(g10784C),.A2(g4467C),.A1(g10727C));
AND2_X1 U_g8174C (.ZN(g8174C),.A2(FE_OFN89_I11360C),.A1(g38C));
AND2_X1 U_g6332C (.ZN(g6332C),.A2(FE_OFN180_g5354C),.A1(g1374C));
AND2_X1 U_g5067C (.ZN(g5067C),.A2(g4811C),.A1(g305C));
AND2_X1 U_g5418C (.ZN(g5418C),.A2(FE_OFN357_g3521C),.A1(g1512C));
AND2_X1 U_g10297C (.ZN(g10297C),.A2(g10001C),.A1(FE_OFN79_g8700C));
AND2_X1 U_g6353C (.ZN(g6353C),.A2(FE_OFN320_g5361C),.A1(g299C));
AND2_X1 U_g11026C (.ZN(g11026C),.A2(FE_OFN14_g10702C),.A1(g386C));
AND2_X1 U_g11212C (.ZN(g11212C),.A2(FE_OFN279_g11157C),.A1(g944C));
AND2_X1 U_g6744C (.ZN(g6744C),.A2(FE_OFN218_g5557C),.A1(g4828C));
AND2_X1 U_g5493C (.ZN(g5493C),.A2(FE_OFN333_g4294C),.A1(g1923C));
AND2_X1 U_g10671C (.ZN(g10671C),.A2(g9473C),.A1(g10411C));
AND2_X1 U_g4383C (.ZN(g4383C),.A2(FE_OFN141_g3829C),.A1(g2517C));
AND2_X1 U_g5256C (.ZN(g5256C),.A2(g627C),.A1(g4297C));
AND2_X1 U_g4220C (.ZN(g4220C),.A2(g3539C),.A1(g105C));
AND2_X1 U_g8380C (.ZN(g8380C),.A2(FE_OFN333_g4294C),.A1(g8252C));
AND2_X1 U_g7071C (.ZN(g7071C),.A2(g6586C),.A1(g5030C));
AND2_X1 U_g4779C (.ZN(g4779C),.A2(FE_OFN307_g4010C),.A1(g501C));
AND2_X1 U_g9613C (.ZN(g9613C),.A2(FE_OFN46_g9125C),.A1(g1176C));
AND2_X1 U_g7705C (.ZN(g7705C),.A2(g4336C),.A1(g5935C));
AND2_X1 U_g9269C (.ZN(g9269C),.A2(FE_OFN266_g18C),.A1(g8933C));
AND2_X1 U_g5181C (.ZN(g5181C),.A2(g802C),.A1(g806C));
AND2_X1 U_g4977C (.ZN(g4977C),.A2(g4807C),.A1(g4567C));
AND2_X1 U_g7948C (.ZN(g7948C),.A2(g7497C),.A1(g70C));
AND2_X1 U_g11149C (.ZN(g11149C),.A2(FE_OFN278_g10927C),.A1(g324C));
AND2_X1 U_g9862C (.ZN(g9862C),.A2(g9778C),.A1(g1601C));
AND2_X1 U_g11387C (.ZN(g11387C),.A2(g3629C),.A1(g11077C));
AND2_X1 U_g7955C (.ZN(g7955C),.A2(g7516C),.A1(g76C));
AND2_X1 U_g4161C (.ZN(g4161C),.A2(g3060C),.A1(FE_OFN251_g1801C));
AND2_X1 U_g11148C (.ZN(g11148C),.A2(g10788C),.A1(g2321C));
AND2_X1 U_g9712C (.ZN(g9712C),.A2(FE_OFN70_g9490C),.A1(g1528C));
AND2_X1 U_g8931C (.ZN(g8931C),.A2(g8164C),.A1(g8642C));
AND2_X1 U_g11097C (.ZN(g11097C),.A2(g10883C),.A1(g378C));
AND3_X1 U_g5421C (.ZN(g5421C),.A3(g3819C),.A2(g109C),.A1(FE_OFN184_I7048C));
AND2_X1 U_g11104C (.ZN(g11104C),.A2(g10937C),.A1(g2963C));
AND2_X1 U_g5263C (.ZN(g5263C),.A2(FE_OFN335_g4737C),.A1(g709C));
AND2_X1 U_g6092C (.ZN(g6092C),.A2(FE_OFN273_g85C),.A1(g1059C));
AND2_X1 U_g4999C (.ZN(g4999C),.A2(FE_OFN154_g4640C),.A1(g1499C));
AND4_X1 U_I6338C (.ZN(I6338C),.A4(g2446C),.A3(g2451C),.A2(g2456C),.A1(g2475C));
AND3_X1 U_g7409C (.ZN(g7409C),.A3(g6858C),.A2(g632C),.A1(g4976C));
AND2_X1 U_g4103C (.ZN(g4103C),.A2(g3060C),.A1(FE_OFN247_g1771C));
AND4_X1 U_I6309C (.ZN(I6309C),.A4(g2475C),.A3(g2456C),.A2(g2451C),.A1(g2446C));
AND2_X1 U_g6580C (.ZN(g6580C),.A2(g5944C),.A1(FE_OFN251_g1801C));
AND2_X1 U_g5631C (.ZN(g5631C),.A2(FE_OFN291_g4880C),.A1(g1056C));
AND2_X1 U_g9414C (.ZN(g9414C),.A2(g9052C),.A1(g1730C));
AND2_X1 U_g9660C (.ZN(g9660C),.A2(FE_OFN45_g9125C),.A1(g1188C));
AND2_X1 U_g9946C (.ZN(g9946C),.A2(FE_OFN68_g9392C),.A1(g9926C));
AND2_X1 U_g5257C (.ZN(g5257C),.A2(FE_OFN335_g4737C),.A1(g691C));
AND2_X1 U_g4732C (.ZN(g4732C),.A2(FE_OFN300_g4002C),.A1(g391C));
AND2_X1 U_g3108C (.ZN(g3108C),.A2(I6331C),.A1(I6330C));
AND2_X1 U_g4753C (.ZN(g4753C),.A2(FE_OFN307_g4010C),.A1(g481C));
AND2_X1 U_g9903C (.ZN(g9903C),.A2(g9673C),.A1(g9885C));
AND2_X1 U_g10625C (.ZN(g10625C),.A2(FE_OFN369_g4525C),.A1(g10454C));
AND2_X1 U_g5605C (.ZN(g5605C),.A2(g704C),.A1(g4828C));
AND2_X1 U_g6623C (.ZN(g6623C),.A2(FE_OFN97_I8869C),.A1(g55C));
AND2_X1 U_g11228C (.ZN(g11228C),.A2(g11060C),.A1(g466C));
AND2_X1 U_g11011C (.ZN(g11011C),.A2(g10809C),.A1(g1968C));
AND2_X1 U_g6889C (.ZN(g6889C),.A2(FE_OFN213_g6003C),.A1(g1941C));
AND2_X1 U_g8040C (.ZN(g8040C),.A2(FE_OFN305_g5151C),.A1(g7523C));
AND2_X1 U_g7822C (.ZN(g7822C),.A2(FE_OFN209_g6863C),.A1(g1914C));
AND2_X1 U_g8123C (.ZN(g8123C),.A2(g7952C),.A1(g1918C));
AND2_X1 U_g11582C (.ZN(g11582C),.A2(g11539C),.A1(g1311C));
AND2_X1 U_g4316C (.ZN(g4316C),.A2(g3275C),.A1(g1965C));
AND2_X1 U_g10969C (.ZN(g10969C),.A2(g10809C),.A1(g3625C));
AND2_X1 U_g5041C (.ZN(g5041C),.A2(FE_OFN223_g4401C),.A1(g3983C));
AND2_X1 U_g9335C (.ZN(g9335C),.A2(FE_OFN275_g48C),.A1(g8975C));
AND2_X1 U_g9831C (.ZN(g9831C),.A2(FE_OFN34_g9785C),.A1(g9727C));
AND2_X1 U_g4565C (.ZN(g4565C),.A2(g4010C),.A1(g534C));
AND2_X1 U_g9422C (.ZN(g9422C),.A2(FE_OFN50_g9030C),.A1(g1750C));
AND2_X1 U_g8648C (.ZN(g8648C),.A2(g8511C),.A1(g4588C));
AND3_X1 U_g8875C (.ZN(g8875C),.A3(g8858C),.A2(FE_OFN92_g2216C),.A1(g8255C));
AND2_X1 U_g5168C (.ZN(g5168C),.A2(g4679C),.A1(g1512C));
AND2_X1 U_g7895C (.ZN(g7895C),.A2(FE_OFN334_g7045C),.A1(g7503C));
AND2_X1 U_g8655C (.ZN(g8655C),.A2(FE_OFN298_g3015C),.A1(g8267C));
AND2_X1 U_g4914C (.ZN(g4914C),.A2(FE_OFN290_g4880C),.A1(g1062C));
AND2_X1 U_g9947C (.ZN(g9947C),.A2(g9392C),.A1(g9927C));
AND2_X1 U_g5772C (.ZN(g5772C),.A2(FE_OFN321_g5261C),.A1(g1555C));
AND2_X1 U_g6838C (.ZN(g6838C),.A2(FE_OFN180_g5354C),.A1(g192C));
AND2_X1 U_g5531C (.ZN(g5531C),.A2(g4290C),.A1(g1666C));
AND2_X1 U_g6795C (.ZN(g6795C),.A2(g5878C),.A1(g5036C));
AND2_X1 U_g10503C (.ZN(g10503C),.A2(FE_OFN336_g1690C),.A1(g9995C));
AND2_X1 U_g8010C (.ZN(g8010C),.A2(g7438C),.A1(g7738C));
AND2_X1 U_g8410C (.ZN(g8410C),.A2(g8146C),.A1(g713C));
AND2_X1 U_g6231C (.ZN(g6231C),.A2(g5608C),.A1(g818C));
AND2_X1 U_g10581C (.ZN(g10581C),.A2(g9473C),.A1(g10336C));
AND2_X1 U_g10450C (.ZN(g10450C),.A2(FE_OFN235_g2024C),.A1(g10364C));
AND2_X1 U_g2804C (.ZN(g2804C),.A2(g1891C),.A1(g2132C));
AND2_X1 U_g3418C (.ZN(g3418C),.A2(FE_OFN352_g109C),.A1(g2379C));
AND2_X1 U_g9653C (.ZN(g9653C),.A2(FE_OFN45_g9125C),.A1(g1185C));
AND2_X1 U_g6205C (.ZN(g6205C),.A2(FE_OFN306_g5128C),.A1(g1515C));
AND2_X1 U_g10818C (.ZN(g10818C),.A2(FE_OFN204_g3664C),.A1(I16220C));
AND2_X1 U_g8172C (.ZN(g8172C),.A2(FE_OFN89_I11360C),.A1(g37C));
AND2_X1 U_g10496C (.ZN(g10496C),.A2(FE_OFN234_g2024C),.A1(g10429C));
AND2_X1 U_g5074C (.ZN(g5074C),.A2(g4608C),.A1(g1771C));
AND2_X1 U_g9869C (.ZN(g9869C),.A2(g9814C),.A1(g1558C));
AND2_X1 U_g9719C (.ZN(g9719C),.A2(g9490C),.A1(g1543C));
AND2_X1 U_g10741C (.ZN(g10741C),.A2(FE_OFN133_g3015C),.A1(g10635C));
AND2_X1 U_g3381C (.ZN(g3381C),.A2(g2756C),.A1(g940C));
AND2_X1 U_g5863C (.ZN(g5863C),.A2(g622C),.A1(g255C));
AND2_X1 U_g8693C (.ZN(g8693C),.A2(g8509C),.A1(g3738C));
AND2_X1 U_g5480C (.ZN(g5480C),.A2(FE_OFN366_g3521C),.A1(g554C));
AND2_X1 U_g4581C (.ZN(g4581C),.A2(g2047C),.A1(g3766C));
AND2_X1 U_g3685C (.ZN(g3685C),.A2(g2981C),.A1(FE_OFN238_g1781C));
AND2_X1 U_g5569C (.ZN(g5569C),.A2(g2338C),.A1(g4816C));
AND2_X1 U_g8555C (.ZN(g8555C),.A2(FE_OFN189_g7638C),.A1(g8409C));
AND2_X1 U_g3263C (.ZN(g3263C),.A2(g2328C),.A1(g2503C));
AND2_X1 U_g9364C (.ZN(g9364C),.A2(g9223C),.A1(g965C));
AND2_X1 U_g4784C (.ZN(g4784C),.A2(FE_OFN307_g4010C),.A1(g506C));
AND2_X4 U_g9454C (.ZN(g9454C),.A2(FE_OFN275_g48C),.A1(g8994C));
AND4_X1 U_I6331C (.ZN(I6331C),.A4(g2077C),.A3(g2074C),.A2(g2070C),.A1(g2060C));
AND2_X1 U_g11299C (.ZN(g11299C),.A2(g11243C),.A1(g4576C));
AND2_X1 U_g6983C (.ZN(g6983C),.A2(FE_OFN343_I5565C),.A1(g6592C));
AND2_X1 U_g7958C (.ZN(g7958C),.A2(FE_OFN198_g7697C),.A1(g736C));
AND2_X1 U_g4995C (.ZN(g4995C),.A2(FE_OFN153_g4640C),.A1(g1474C));
AND2_X1 U_g4079C (.ZN(g4079C),.A2(g2276C),.A1(FE_OFN237_g1806C));
AND2_X1 U_g2264C (.ZN(g2264C),.A2(g1766C),.A1(FE_OFN247_g1771C));
AND2_X1 U_g2160C (.ZN(g2160C),.A2(g746C),.A1(g745C));
AND2_X1 U_g3257C (.ZN(g3257C),.A2(g2496C),.A1(g378C));
AND2_X1 U_g3101C (.ZN(g3101C),.A2(I6310C),.A1(I6309C));
AND2_X1 U_g5000C (.ZN(g5000C),.A2(FE_OFN153_g4640C),.A1(g1470C));
AND2_X1 U_g3301C (.ZN(g3301C),.A2(g2544C),.A1(g1346C));
AND2_X1 U_g5126C (.ZN(g5126C),.A2(g4671C),.A1(g1104C));
AND4_X1 U_I5084C (.ZN(I5084C),.A4(g1478C),.A3(g1474C),.A2(g1470C),.A1(g1462C));
AND2_X1 U_g9412C (.ZN(g9412C),.A2(g9052C),.A1(g1727C));
AND2_X1 U_g9389C (.ZN(g9389C),.A2(FE_OFN47_g9151C),.A1(g1330C));
AND2_X1 U_g2379C (.ZN(g2379C),.A2(g743C),.A1(g744C));
AND2_X1 U_g10706C (.ZN(g10706C),.A2(FE_OFN345_g3015C),.A1(g10567C));
AND3_X1 U_I16145C (.ZN(I16145C),.A3(g10446C),.A2(g10447C),.A1(g10366C));
AND2_X1 U_g10597C (.ZN(g10597C),.A2(FE_OFN369_g4525C),.A1(g10533C));
AND3_X1 U_g8965C (.ZN(g8965C),.A3(g8849C),.A2(FE_OFN281_g2216C),.A1(g8110C));
AND2_X1 U_g5608C (.ZN(g5608C),.A2(g4831C),.A1(g814C));
AND2_X1 U_g5220C (.ZN(g5220C),.A2(g4776C),.A1(g1083C));
AND2_X1 U_g10624C (.ZN(g10624C),.A2(FE_OFN370_g4525C),.A1(g10494C));
AND2_X1 U_g10300C (.ZN(g10300C),.A2(g10019C),.A1(FE_OFN76_g8700C));
AND2_X1 U_g5023C (.ZN(g5023C),.A2(FE_OFN288_g4263C),.A1(g1071C));
AND2_X1 U_g4432C (.ZN(g4432C),.A2(g1975C),.A1(g3723C));
AND2_X1 U_g4053C (.ZN(g4053C),.A2(FE_OFN224_g2276C),.A1(FE_OFN253_g1786C));
AND2_X1 U_g8050C (.ZN(g8050C),.A2(FE_OFN177_g5919C),.A1(g7596C));
AND2_X1 U_g5588C (.ZN(g5588C),.A2(FE_OFN367_g3521C),.A1(g1639C));
AND3_X1 U_g6679C (.ZN(g6679C),.A3(g109C),.A2(g6074C),.A1(FE_OFN184_I7048C));
AND2_X1 U_g9963C (.ZN(g9963C),.A2(FE_OFN280_g9536C),.A1(g9953C));
AND2_X1 U_g3772C (.ZN(g3772C),.A2(g3089C),.A1(g2542C));
AND2_X1 U_g5051C (.ZN(g5051C),.A2(g2506C),.A1(g4432C));
AND2_X1 U_g6831C (.ZN(g6831C),.A2(FE_OFN179_g5354C),.A1(g207C));
AND2_X1 U_g2981C (.ZN(g2981C),.A2(g2264C),.A1(FE_OFN236_g1776C));
AND2_X1 U_g8724C (.ZN(g8724C),.A2(g7910C),.A1(g8214C));
AND2_X1 U_g4157C (.ZN(g4157C),.A2(g3060C),.A1(FE_OFN239_g1796C));
AND2_X1 U_g9707C (.ZN(g9707C),.A2(g9474C),.A1(g1583C));
AND3_X1 U_g8878C (.ZN(g8878C),.A3(FE_OFN73_g8858C),.A2(FE_OFN93_g2216C),.A1(g8099C));
AND2_X1 U_g2132C (.ZN(g2132C),.A2(g1882C),.A1(g1872C));
AND2_X1 U_g10763C (.ZN(g10763C),.A2(FE_OFN345_g3015C),.A1(g10639C));
AND3_X1 U_g8289C (.ZN(g8289C),.A3(g2216C),.A2(g8109C),.A1(g6777C));
AND2_X1 U_g7898C (.ZN(g7898C),.A2(g7045C),.A1(g7511C));
AND2_X1 U_g11271C (.ZN(g11271C),.A2(g11203C),.A1(g4753C));
AND2_X1 U_g11461C (.ZN(g11461C),.A2(FE_OFN100_g4421C),.A1(g11225C));
AND2_X1 U_g5732C (.ZN(g5732C),.A2(FE_OFN353_g5117C),.A1(g1604C));
AND2_X1 U_g11145C (.ZN(g11145C),.A2(FE_OFN278_g10927C),.A1(g315C));
AND2_X1 U_g11031C (.ZN(g11031C),.A2(FE_OFN14_g10702C),.A1(g411C));
AND2_X1 U_g9865C (.ZN(g9865C),.A2(g9773C),.A1(g1607C));
AND2_X1 U_g5944C (.ZN(g5944C),.A2(g5233C),.A1(g1796C));
AND2_X1 U_g9715C (.ZN(g9715C),.A2(FE_OFN70_g9490C),.A1(g1531C));
AND2_X1 U_g9604C (.ZN(g9604C),.A2(FE_OFN51_g9111C),.A1(g1194C));
AND2_X1 U_g8799C (.ZN(g8799C),.A2(FE_OFN331_g8696C),.A1(g8647C));
AND2_X1 U_g11198C (.ZN(g11198C),.A2(FE_OFN15_g10702C),.A1(g4778C));
AND2_X1 U_g6873C (.ZN(g6873C),.A2(g6557C),.A1(g3263C));
AND2_X1 U_g6632C (.ZN(g6632C),.A2(FE_OFN283_I8869C),.A1(g61C));
AND2_X1 U_g6095C (.ZN(g6095C),.A2(FE_OFN273_g85C),.A1(g1062C));
AND2_X1 U_g3863C (.ZN(g3863C),.A2(g1696C),.A1(g1703C));
AND2_X1 U_g9833C (.ZN(g9833C),.A2(FE_OFN34_g9785C),.A1(g9729C));
AND2_X1 U_g6653C (.ZN(g6653C),.A2(I8869C),.A1(g70C));
AND2_X1 U_g6102C (.ZN(g6102C),.A2(FE_OFN273_g85C),.A1(g1038C));
AND2_X1 U_g7819C (.ZN(g7819C),.A2(FE_OFN206_g6863C),.A1(g1887C));
AND2_X1 U_g11393C (.ZN(g11393C),.A2(g7914C),.A1(g11280C));
AND2_X1 U_g2511C (.ZN(g2511C),.A2(g456C),.A1(FE_OFN254_g461C));
AND2_X1 U_g7088C (.ZN(g7088C),.A2(g6432C),.A1(g2331C));
AND2_X1 U_g9584C (.ZN(g9584C),.A2(FE_OFN53_g9173C),.A1(g1341C));
AND2_X1 U_g9896C (.ZN(g9896C),.A2(FE_OFN60_g9624C),.A1(g9696C));
AND3_X1 U_g8209C (.ZN(g8209C),.A3(g7622C),.A2(g3068C),.A1(g4094C));
AND2_X1 U_g6752C (.ZN(g6752C),.A2(g2343C),.A1(g6187C));
AND2_X1 U_g4778C (.ZN(g4778C),.A2(g4002C),.A1(g421C));
AND2_X1 U_g11161C (.ZN(g11161C),.A2(g10937C),.A1(g1969C));
AND2_X1 U_g9268C (.ZN(g9268C),.A2(g8947C),.A1(g6109C));
AND2_X1 U_g5681C (.ZN(g5681C),.A2(FE_OFN365_g5361C),.A1(g135C));
AND2_X1 U_g7951C (.ZN(g7951C),.A2(g7505C),.A1(g73C));
AND2_X1 U_g9419C (.ZN(g9419C),.A2(FE_OFN50_g9030C),.A1(g1744C));
AND2_X1 U_g10268C (.ZN(g10268C),.A2(FE_OFN267_g109C),.A1(I15287C));
AND2_X1 U_g5533C (.ZN(g5533C),.A2(g4292C),.A1(g1724C));
AND2_X4 U_g9052C (.ZN(g9052C),.A2(FE_OFN276_g48C),.A1(g8936C));
AND2_X1 U_g6786C (.ZN(g6786C),.A2(g5919C),.A1(g178C));
AND2_X1 U_g10670C (.ZN(g10670C),.A2(g9097C),.A1(g10396C));
AND2_X1 U_g11087C (.ZN(g11087C),.A2(FE_OFN4_g10950C),.A1(g829C));
AND2_X1 U_g4949C (.ZN(g4949C),.A2(g4449C),.A1(I5815C));
AND2_X1 U_g6364C (.ZN(g6364C),.A2(FE_OFN346_g4381C),.A1(g5851C));
AND2_X1 U_g7825C (.ZN(g7825C),.A2(FE_OFN206_g6863C),.A1(g1941C));
AND2_X1 U_g4998C (.ZN(g4998C),.A2(FE_OFN303_g4678C),.A1(g1304C));
AND2_X1 U_g10667C (.ZN(g10667C),.A2(g9424C),.A1(g10405C));
AND2_X1 U_g7136C (.ZN(g7136C),.A2(g6718C),.A1(g5190C));
AND2_X1 U_g6532C (.ZN(g6532C),.A2(FE_OFN282_g6165C),.A1(g339C));
AND2_X1 U_g9385C (.ZN(g9385C),.A2(FE_OFN48_g9151C),.A1(g1324C));
AND4_X1 U_I5690C (.ZN(I5690C),.A4(g1448C),.A3(g1444C),.A2(g1440C),.A1(g1436C));
AND2_X1 U_g4484C (.ZN(g4484C),.A2(FE_OFN302_g3913C),.A1(g1137C));
AND2_X1 U_g9897C (.ZN(g9897C),.A2(FE_OFN60_g9624C),.A1(g9699C));
AND2_X1 U_g9425C (.ZN(g9425C),.A2(FE_OFN49_g9030C),.A1(g1753C));
AND2_X1 U_g3383C (.ZN(g3383C),.A2(FE_OFN324_g18C),.A1(g186C));
AND2_X1 U_g5601C (.ZN(g5601C),.A2(g4880C),.A1(g1035C));
AND2_X1 U_g7943C (.ZN(g7943C),.A2(g7467C),.A1(g64C));
AND2_X1 U_g11171C (.ZN(g11171C),.A2(FE_OFN21_g10702C),.A1(g481C));
AND2_X1 U_g3423C (.ZN(g3423C),.A2(I6631C),.A1(I6630C));
AND2_X1 U_g7230C (.ZN(g7230C),.A2(g6447C),.A1(g6064C));
AND2_X1 U_g4952C (.ZN(g4952C),.A2(FE_OFN299_g4457C),.A1(g1648C));
AND2_X1 U_g6787C (.ZN(g6787C),.A2(FE_OFN319_g5361C),.A1(g266C));
AND3_X1 U_g8968C (.ZN(g8968C),.A3(g8849C),.A2(FE_OFN281_g2216C),.A1(g8089C));
AND2_X1 U_g10306C (.ZN(g10306C),.A2(g9082C),.A1(g10007C));
AND2_X1 U_g9331C (.ZN(g9331C),.A2(FE_OFN275_g48C),.A1(g8972C));
AND2_X1 U_g11459C (.ZN(g11459C),.A2(FE_OFN100_g4421C),.A1(g11221C));
AND2_X1 U_g4561C (.ZN(g4561C),.A2(g4010C),.A1(g538C));
AND2_X1 U_g11425C (.ZN(g11425C),.A2(g10629C),.A1(I16982C));
AND2_X1 U_g11458C (.ZN(g11458C),.A2(FE_OFN99_g4421C),.A1(g11219C));
AND2_X1 U_g5739C (.ZN(g5739C),.A2(FE_OFN315_g5117C),.A1(g1607C));
AND2_X1 U_g7496C (.ZN(g7496C),.A2(g64C),.A1(FE_OFN83_g2176C));
AND2_X1 U_g4986C (.ZN(g4986C),.A2(FE_OFN146_g4682C),.A1(g1411C));
AND2_X1 U_g11010C (.ZN(g11010C),.A2(FE_OFN18_g10702C),.A1(g5187C));
AND2_X1 U_g3999C (.ZN(g3999C),.A2(g2777C),.A1(g1741C));
AND2_X1 U_g8175C (.ZN(g8175C),.A2(FE_OFN89_I11360C),.A1(g39C));
AND2_X1 U_g8722C (.ZN(g8722C),.A2(g7908C),.A1(g8210C));
AND2_X1 U_g4764C (.ZN(g4764C),.A2(FE_OFN300_g4002C),.A1(g411C));
AND2_X1 U_g7137C (.ZN(g7137C),.A2(g6354C),.A1(g5590C));
AND2_X1 U_g7891C (.ZN(g7891C),.A2(FE_OFN334_g7045C),.A1(g7471C));
AND2_X1 U_g8651C (.ZN(g8651C),.A2(FE_OFN348_g3015C),.A1(g8261C));
AND2_X1 U_g5479C (.ZN(g5479C),.A2(g4243C),.A1(g1845C));
AND2_X1 U_g11599C (.ZN(g11599C),.A2(g11575C),.A1(g1341C));
AND2_X1 U_g6684C (.ZN(g6684C),.A2(g5836C),.A1(g91C));
AND2_X1 U_g6745C (.ZN(g6745C),.A2(FE_OFN218_g5557C),.A1(g5605C));
AND2_X1 U_g6639C (.ZN(g6639C),.A2(FE_OFN282_g6165C),.A1(g357C));
AND2_X1 U_g10937C (.ZN(g10937C),.A2(FE_OFN13_g10702C),.A1(g4822C));
AND2_X1 U_g3696C (.ZN(g3696C),.A2(FE_OFN364_g3015C),.A1(g1713C));
AND2_X1 U_g4503C (.ZN(g4503C),.A2(g3943C),.A1(g654C));
AND2_X1 U_g6791C (.ZN(g6791C),.A2(FE_OFN319_g5361C),.A1(g269C));
AND2_X1 U_g5190C (.ZN(g5190C),.A2(g4678C),.A1(g1245C));
AND2_X1 U_g5390C (.ZN(g5390C),.A2(g4671C),.A1(g1101C));
AND2_X1 U_g8384C (.ZN(g8384C),.A2(FE_OFN325_g18C),.A1(g8180C));
AND2_X1 U_g4224C (.ZN(g4224C),.A2(FE_OFN132_g3015C),.A1(g1092C));
AND2_X1 U_g5501C (.ZN(g5501C),.A2(g4273C),.A1(g1672C));
AND2_X4 U_g9173C (.ZN(g9173C),.A2(FE_OFN276_g48C),.A1(g8968C));
AND2_X1 U_g6759C (.ZN(g6759C),.A2(g5919C),.A1(g148C));
AND2_X1 U_g8838C (.ZN(g8838C),.A2(FE_OFN328_g8709C),.A1(g8602C));
AND2_X1 U_g8024C (.ZN(g8024C),.A2(FE_OFN322_g4449C),.A1(g6577C));
AND2_X1 U_g10666C (.ZN(g10666C),.A2(g9424C),.A1(g10402C));
AND2_X1 U_g11158C (.ZN(g11158C),.A2(FE_OFN278_g10927C),.A1(g309C));
AND2_X1 U_g9602C (.ZN(g9602C),.A2(g9010C),.A1(g932C));
AND2_X1 U_g5704C (.ZN(g5704C),.A2(FE_OFN164_g5361C),.A1(g143C));
AND2_X1 U_g4617C (.ZN(g4617C),.A2(g3879C),.A1(g3275C));
AND2_X2 U_g11561C (.ZN(g11561C),.A2(FE_OFN364_g3015C),.A1(g11492C));
AND2_X1 U_g9868C (.ZN(g9868C),.A2(g9814C),.A1(g1555C));
AND2_X1 U_g11295C (.ZN(g11295C),.A2(g11239C),.A1(g4554C));
AND2_X1 U_g11144C (.ZN(g11144C),.A2(FE_OFN10_g10702C),.A1(g305C));
AND2_X1 U_g9718C (.ZN(g9718C),.A2(FE_OFN70_g9490C),.A1(g1540C));
AND2_X1 U_g3434C (.ZN(g3434C),.A2(g2355C),.A1(g237C));
AND2_X1 U_g4987C (.ZN(g4987C),.A2(FE_OFN147_g4682C),.A1(g1440C));
AND2_X1 U_g4771C (.ZN(g4771C),.A2(FE_OFN307_g4010C),.A1(g496C));
AND2_X1 U_g5250C (.ZN(g5250C),.A2(g4678C),.A1(g1270C));
AND2_X1 U_g6098C (.ZN(g6098C),.A2(FE_OFN273_g85C),.A1(g1065C));
AND2_X1 U_g9582C (.ZN(g9582C),.A2(FE_OFN53_g9173C),.A1(g2725C));
AND2_X1 U_g6833C (.ZN(g6833C),.A2(FE_OFN178_g5354C),.A1(g186C));
AND2_X1 U_g3533C (.ZN(g3533C),.A2(g2892C),.A1(g1981C));
AND2_X1 U_g4892C (.ZN(g4892C),.A2(g4739C),.A1(g632C));
AND2_X1 U_g8104C (.ZN(g8104C),.A2(g7852C),.A1(g5493C));
AND2_X1 U_g9415C (.ZN(g9415C),.A2(FE_OFN54_g9052C),.A1(g1733C));
AND2_X1 U_g8499C (.ZN(g8499C),.A2(g4737C),.A1(g8377C));
AND2_X1 U_g9664C (.ZN(g9664C),.A2(FE_OFN46_g9125C),.A1(g1191C));
AND2_X1 U_g9721C (.ZN(g9721C),.A2(FE_OFN359_g18C),.A1(g9413C));
AND2_X1 U_g6162C (.ZN(g6162C),.A2(g5200C),.A1(g3584C));
AND2_X1 U_g4991C (.ZN(g4991C),.A2(FE_OFN154_g4640C),.A1(g1508C));
AND2_X1 U_g6362C (.ZN(g6362C),.A2(FE_OFN346_g4381C),.A1(g5846C));
AND4_X1 U_I6631C (.ZN(I6631C),.A4(FE_OFN237_g1806C),.A3(FE_OFN251_g1801C),.A2(FE_OFN239_g1796C),.A1(FE_OFN252_g1791C));
AND2_X1 U_g10685C (.ZN(g10685C),.A2(FE_OFN136_g3863C),.A1(g10383C));
AND2_X1 U_g4340C (.ZN(g4340C),.A2(FE_OFN351_g3913C),.A1(g1153C));
AND2_X1 U_g11023C (.ZN(g11023C),.A2(g10702C),.A1(g440C));
AND2_X1 U_g8044C (.ZN(g8044C),.A2(FE_OFN177_g5919C),.A1(g7598C));
AND2_X1 U_g11224C (.ZN(g11224C),.A2(g11157C),.A1(g968C));
AND2_X1 U_g11571C (.ZN(g11571C),.A2(g11561C),.A1(g2018C));
AND2_X1 U_g4959C (.ZN(g4959C),.A2(FE_OFN147_g4682C),.A1(g1520C));
AND2_X1 U_g10334C (.ZN(g10334C),.A2(FE_OFN267_g109C),.A1(I15365C));
AND2_X1 U_g5626C (.ZN(g5626C),.A2(FE_OFN367_g3521C),.A1(g1633C));
AND2_X1 U_g9940C (.ZN(g9940C),.A2(FE_OFN67_g9367C),.A1(g9920C));
AND2_X1 U_g4876C (.ZN(g4876C),.A2(FE_OFN132_g3015C),.A1(g1086C));
AND2_X1 U_g6728C (.ZN(g6728C),.A2(FE_OFN310_g4336C),.A1(g4482C));
AND2_X1 U_g6730C (.ZN(g6730C),.A2(g5013C),.A1(g1872C));
AND2_X1 U_g9689C (.ZN(g9689C),.A2(FE_OFN59_g9432C),.A1(g263C));
AND2_X1 U_g10762C (.ZN(g10762C),.A2(FE_OFN131_g3015C),.A1(g10635C));
AND2_X1 U_g6070C (.ZN(g6070C),.A2(FE_OFN273_g85C),.A1(g1050C));
AND2_X1 U_g9428C (.ZN(g9428C),.A2(FE_OFN50_g9030C),.A1(g1756C));
AND2_X4 U_g9030C (.ZN(g9030C),.A2(FE_OFN276_g48C),.A1(g8935C));
AND2_X1 U_g9430C (.ZN(g9430C),.A2(FE_OFN49_g9030C),.A1(g1759C));
AND2_X1 U_g8927C (.ZN(g8927C),.A2(g8642C),.A1(g2216C));
AND2_X1 U_g7068C (.ZN(g7068C),.A2(g6586C),.A1(g5024C));
AND2_X1 U_g8014C (.ZN(g8014C),.A2(g7438C),.A1(g7740C));
AND2_X1 U_g11392C (.ZN(g11392C),.A2(g7914C),.A1(g11278C));
AND2_X1 U_g5782C (.ZN(g5782C),.A2(g5222C),.A1(g1558C));
AND2_X1 U_g4824C (.ZN(g4824C),.A2(g4099C),.A1(g774C));
AND2_X1 U_g6331C (.ZN(g6331C),.A2(FE_OFN180_g5354C),.A1(g201C));
AND2_X1 U_g4236C (.ZN(g4236C),.A2(FE_OFN132_g3015C),.A1(g1098C));
AND2_X1 U_g11559C (.ZN(g11559C),.A2(FE_OFN27_g11519C),.A1(FE_OFN251_g1801C));
AND2_X1 U_g9609C (.ZN(g9609C),.A2(FE_OFN42_g9205C),.A1(g907C));
AND2_X1 U_g11558C (.ZN(g11558C),.A2(FE_OFN27_g11519C),.A1(FE_OFN239_g1796C));
AND2_X1 U_g6087C (.ZN(g6087C),.A2(FE_OFN271_g85C),.A1(g1056C));
AND2_X1 U_g5526C (.ZN(g5526C),.A2(g4294C),.A1(g1950C));
AND2_X1 U_g10751C (.ZN(g10751C),.A2(FE_OFN133_g3015C),.A1(g10646C));
AND2_X1 U_g10772C (.ZN(g10772C),.A2(FE_OFN345_g3015C),.A1(g10655C));
AND2_X1 U_g8135C (.ZN(g8135C),.A2(g7883C),.A1(g1945C));
AND2_X1 U_g11544C (.ZN(g11544C),.A2(g10584C),.A1(g11515C));
AND2_X1 U_g5084C (.ZN(g5084C),.A2(FE_OFN299_g4457C),.A1(g1776C));
AND2_X1 U_g8382C (.ZN(g8382C),.A2(FE_OFN196_g7697C),.A1(g5248C));
AND2_X1 U_g10230C (.ZN(g10230C),.A2(g9968C),.A1(g8700C));
AND2_X1 U_g5484C (.ZN(g5484C),.A2(FE_OFN333_g4294C),.A1(g1896C));
AND2_X1 U_g7241C (.ZN(g7241C),.A2(g5557C),.A1(g6772C));
AND2_X1 U_g3942C (.ZN(g3942C),.A2(FE_OFN260_g18C),.A1(g219C));
AND2_X1 U_g10638C (.ZN(g10638C),.A2(g3829C),.A1(g10383C));
AND2_X1 U_g4064C (.ZN(g4064C),.A2(g2774C),.A1(g1759C));
AND2_X1 U_g9365C (.ZN(g9365C),.A2(FE_OFN48_g9151C),.A1(g1321C));
AND2_X1 U_g9861C (.ZN(g9861C),.A2(g9579C),.A1(g9738C));
AND2_X1 U_g11255C (.ZN(g11255C),.A2(g11060C),.A1(g456C));
AND2_X1 U_g11189C (.ZN(g11189C),.A2(FE_OFN15_g10702C),.A1(g4736C));
AND2_X1 U_g10510C (.ZN(g10510C),.A2(FE_OFN336_g1690C),.A1(g10019C));
AND3_X1 U_g8947C (.ZN(g8947C),.A3(g8828C),.A2(FE_OFN92_g2216C),.A1(g8056C));
AND2_X1 U_g2917C (.ZN(g2917C),.A2(g1657C),.A1(g2424C));
AND2_X2 U_g5919C (.ZN(g5919C),.A2(FE_OFN269_g109C),.A1(I7048C));
AND2_X1 U_g11188C (.ZN(g11188C),.A2(FE_OFN15_g10702C),.A1(g4732C));
AND2_X1 U_g9846C (.ZN(g9846C),.A2(g9764C),.A1(g287C));
AND2_X1 U_g7818C (.ZN(g7818C),.A2(FE_OFN206_g6863C),.A1(g1878C));
AND2_X1 U_g11460C (.ZN(g11460C),.A2(FE_OFN99_g4421C),.A1(g11223C));
AND2_X1 U_g5276C (.ZN(g5276C),.A2(FE_OFN335_g4737C),.A1(g736C));
AND2_X1 U_g11030C (.ZN(g11030C),.A2(FE_OFN17_g10702C),.A1(g406C));
AND2_X1 U_g11093C (.ZN(g11093C),.A2(FE_OFN4_g10950C),.A1(g841C));
AND2_X1 U_g7893C (.ZN(g7893C),.A2(FE_OFN334_g7045C),.A1(g7478C));
AND2_X1 U_g8653C (.ZN(g8653C),.A2(FE_OFN348_g3015C),.A1(g8265C));
AND2_X1 U_g10442C (.ZN(g10442C),.A2(FE_OFN245_g1690C),.A1(g9968C));
AND2_X1 U_g6535C (.ZN(g6535C),.A2(g6165C),.A1(g345C));
AND2_X1 U_g8102C (.ZN(g8102C),.A2(g7852C),.A1(g5485C));
AND4_X1 U_I5085C (.ZN(I5085C),.A4(g1508C),.A3(g1504C),.A2(g1494C),.A1(g1490C));
AND2_X1 U_g5004C (.ZN(g5004C),.A2(FE_OFN303_g4678C),.A1(g1296C));
AND2_X1 U_g3912C (.ZN(g3912C),.A2(FE_OFN359_g18C),.A1(g207C));
AND2_X1 U_g7186C (.ZN(g7186C),.A2(g6403C),.A1(g2503C));
AND2_X1 U_g4489C (.ZN(g4489C),.A2(FE_OFN103_g3586C),.A1(g348C));
AND2_X1 U_g9662C (.ZN(g9662C),.A2(g9292C),.A1(g123C));
AND2_X1 U_g9418C (.ZN(g9418C),.A2(FE_OFN56_g9052C),.A1(g1741C));
AND2_X1 U_g11218C (.ZN(g11218C),.A2(FE_OFN279_g11157C),.A1(g959C));
AND2_X1 U_g4471C (.ZN(g4471C),.A2(FE_OFN302_g3913C),.A1(g1121C));
AND2_X1 U_g10746C (.ZN(g10746C),.A2(FE_OFN364_g3015C),.A1(g10643C));
AND2_X1 U_g7125C (.ZN(g7125C),.A2(g5763C),.A1(g1212C));
AND2_X1 U_g7821C (.ZN(g7821C),.A2(FE_OFN209_g6863C),.A1(g1905C));
AND2_X1 U_g6246C (.ZN(g6246C),.A2(FE_OFN164_g5361C),.A1(g178C));
AND2_X1 U_g9256C (.ZN(g9256C),.A2(g8963C),.A1(g6109C));
AND2_X1 U_g8042C (.ZN(g8042C),.A2(FE_OFN305_g5151C),.A1(g7533C));
AND2_X1 U_g10237C (.ZN(g10237C),.A2(g9082C),.A1(g9968C));
AND2_X1 U_g7939C (.ZN(g7939C),.A2(g7460C),.A1(g61C));
AND2_X1 U_g8786C (.ZN(g8786C),.A2(FE_OFN331_g8696C),.A1(g8638C));
AND2_X1 U_g10684C (.ZN(g10684C),.A2(FE_OFN136_g3863C),.A1(g10382C));
AND2_X1 U_g11455C (.ZN(g11455C),.A2(FE_OFN99_g4421C),.A1(g11233C));
AND2_X1 U_g8364C (.ZN(g8364C),.A2(g8146C),.A1(g658C));
AND3_X1 U_g2990C (.ZN(g2990C),.A3(g1814C),.A2(g2557C),.A1(g2061C));
AND2_X1 U_g9847C (.ZN(g9847C),.A2(FE_OFN57_g9432C),.A1(g290C));
AND2_X1 U_g8054C (.ZN(g8054C),.A2(FE_OFN177_g5919C),.A1(g7584C));
AND2_X1 U_g5617C (.ZN(g5617C),.A2(FE_OFN290_g4880C),.A1(g1050C));
AND2_X1 U_g6502C (.ZN(g6502C),.A2(FE_OFN363_I5565C),.A1(g5981C));
AND2_X1 U_g5789C (.ZN(g5789C),.A2(FE_OFN321_g5261C),.A1(g1561C));
AND2_X1 U_g4009C (.ZN(g4009C),.A2(g2774C),.A1(g1747C));
AND2_X1 U_g11277C (.ZN(g11277C),.A2(g11199C),.A1(g4779C));
AND2_X1 U_g6940C (.ZN(g6940C),.A2(g1945C),.A1(g6472C));
AND2_X1 U_g7061C (.ZN(g7061C),.A2(g6760C),.A1(g790C));
AND2_X1 U_g11595C (.ZN(g11595C),.A2(g11575C),.A1(g1336C));
AND2_X1 U_g5771C (.ZN(g5771C),.A2(FE_OFN321_g5261C),.A1(g1534C));
AND2_X1 U_g8553C (.ZN(g8553C),.A2(FE_OFN330_g7638C),.A1(g8405C));
AND2_X1 U_g4836C (.ZN(g4836C),.A2(g3943C),.A1(g643C));
AND2_X1 U_g5547C (.ZN(g5547C),.A2(g4292C),.A1(g1733C));
AND2_X1 U_g6216C (.ZN(g6216C),.A2(FE_OFN306_g5128C),.A1(g1407C));
AND2_X1 U_g4967C (.ZN(g4967C),.A2(FE_OFN146_g4682C),.A1(g1515C));
AND2_X1 U_g6671C (.ZN(g6671C),.A2(FE_OFN282_g6165C),.A1(g342C));
AND2_X1 U_g7200C (.ZN(g7200C),.A2(g6447C),.A1(g3098C));
AND2_X1 U_g3661C (.ZN(g3661C),.A2(g3257C),.A1(g382C));
AND2_X1 U_g7046C (.ZN(g7046C),.A2(g6702C),.A1(g4998C));
AND2_X1 U_g4229C (.ZN(g4229C),.A2(g4673C),.A1(g999C));
AND2_X1 U_g8389C (.ZN(g8389C),.A2(g8220C),.A1(g5263C));
AND2_X1 U_g6430C (.ZN(g6430C),.A2(FE_OFN217_g5013C),.A1(g5044C));
AND2_X1 U_g4993C (.ZN(g4993C),.A2(FE_OFN147_g4682C),.A1(g1448C));
AND2_X1 U_g6247C (.ZN(g6247C),.A2(FE_OFN365_g5361C),.A1(g127C));
AND2_X1 U_g9257C (.ZN(g9257C),.A2(g8964C),.A1(g6109C));
AND2_X1 U_g11170C (.ZN(g11170C),.A2(FE_OFN8_g10702C),.A1(g525C));
AND2_X1 U_g7145C (.ZN(g7145C),.A2(g6718C),.A1(g5250C));
AND2_X1 U_g5738C (.ZN(g5738C),.A2(FE_OFN353_g5117C),.A1(g1586C));
AND2_X1 U_g6826C (.ZN(g6826C),.A2(g5354C),.A1(g225C));
AND2_X1 U_g7191C (.ZN(g7191C),.A2(FE_OFN310_g4336C),.A1(g5219C));
AND2_X1 U_g3998C (.ZN(g3998C),.A2(g2276C),.A1(g2677C));
AND2_X1 U_g6741C (.ZN(g6741C),.A2(FE_OFN219_g5557C),.A1(g3284C));
AND2_X1 U_g5478C (.ZN(g5478C),.A2(FE_OFN333_g4294C),.A1(g1905C));
AND2_X1 U_g11167C (.ZN(g11167C),.A2(FE_OFN8_g10702C),.A1(g538C));
AND2_X1 U_g11194C (.ZN(g11194C),.A2(g10927C),.A1(g4764C));
AND2_X1 U_g11589C (.ZN(g11589C),.A2(g11539C),.A1(g1333C));
AND2_X1 U_g6638C (.ZN(g6638C),.A2(FE_OFN283_I8869C),.A1(g64C));
AND2_X2 U_g4921C (.ZN(g4921C),.A2(g4431C),.A1(g627C));
AND2_X1 U_g7536C (.ZN(g7536C),.A2(g76C),.A1(FE_OFN83_g2176C));
AND2_X1 U_g9585C (.ZN(g9585C),.A2(g8995C),.A1(g889C));
AND2_X1 U_g2957C (.ZN(g2957C),.A2(g1663C),.A1(g2424C));
AND2_X1 U_g11588C (.ZN(g11588C),.A2(g11547C),.A1(g1330C));
AND2_X1 U_g5690C (.ZN(g5690C),.A2(FE_OFN353_g5117C),.A1(g1567C));
AND2_X1 U_g6883C (.ZN(g6883C),.A2(FE_OFN213_g6003C),.A1(g1923C));
AND2_X1 U_g4837C (.ZN(g4837C),.A2(FE_OFN297_g3015C),.A1(g1068C));
AND3_X1 U_g8963C (.ZN(g8963C),.A3(g8849C),.A2(FE_OFN92_g2216C),.A1(g8056C));
AND2_X1 U_g8791C (.ZN(g8791C),.A2(FE_OFN331_g8696C),.A1(g8641C));
AND2_X1 U_g6217C (.ZN(g6217C),.A2(FE_OFN291_g4880C),.A1(g563C));
AND4_X1 U_I6316C (.ZN(I6316C),.A4(g2395C),.A3(g2381C),.A2(g2087C),.A1(g2082C));
AND2_X1 U_g11022C (.ZN(g11022C),.A2(g10702C),.A1(g444C));
AND2_X1 U_g5915C (.ZN(g5915C),.A2(g4977C),.A1(g4168C));
AND2_X1 U_g4788C (.ZN(g4788C),.A2(FE_OFN307_g4010C),.A1(g511C));
AND2_X1 U_g5110C (.ZN(g5110C),.A2(FE_OFN299_g4457C),.A1(FE_OFN237_g1806C));
AND2_X1 U_g11254C (.ZN(g11254C),.A2(g11083C),.A1(g986C));
AND2_X1 U_g6827C (.ZN(g6827C),.A2(FE_OFN178_g5354C),.A1(g219C));
AND3_X1 U_g8957C (.ZN(g8957C),.A3(g8828C),.A2(FE_OFN281_g2216C),.A1(g8081C));
AND2_X1 U_g6333C (.ZN(g6333C),.A2(FE_OFN180_g5354C),.A1(g197C));
AND2_X1 U_g8049C (.ZN(g8049C),.A2(FE_OFN177_g5919C),.A1(g7567C));
AND2_X1 U_g4392C (.ZN(g4392C),.A2(FE_OFN137_g3829C),.A1(g3273C));
AND2_X1 U_g9856C (.ZN(g9856C),.A2(g9773C),.A1(g1592C));
AND2_X1 U_g9411C (.ZN(g9411C),.A2(g9052C),.A1(g1724C));
AND2_X1 U_g5002C (.ZN(g5002C),.A2(FE_OFN154_g4640C),.A1(g1494C));
AND2_X1 U_g11101C (.ZN(g11101C),.A2(FE_OFN4_g10950C),.A1(g857C));
AND2_X1 U_g11177C (.ZN(g11177C),.A2(FE_OFN20_g10702C),.A1(g511C));
AND2_X1 U_g11560C (.ZN(g11560C),.A2(FE_OFN27_g11519C),.A1(g1806C));
AND2_X1 U_g8098C (.ZN(g8098C),.A2(g7852C),.A1(g5478C));
AND2_X1 U_g3970C (.ZN(g3970C),.A2(FE_OFN260_g18C),.A1(g225C));
AND2_X1 U_g4941C (.ZN(g4941C),.A2(FE_OFN290_g4880C),.A1(g1038C));
AND2_X1 U_g10453C (.ZN(g10453C),.A2(FE_OFN234_g2024C),.A1(g10437C));
AND2_X1 U_g5877C (.ZN(g5877C),.A2(g639C),.A1(g4921C));
AND2_X1 U_g6662C (.ZN(g6662C),.A2(FE_OFN282_g6165C),.A1(g366C));
AND2_X1 U_g7935C (.ZN(g7935C),.A2(g7454C),.A1(g58C));
AND2_X1 U_g6067C (.ZN(g6067C),.A2(g85C),.A1(g1047C));
AND4_X1 U_I6317C (.ZN(I6317C),.A4(g2438C),.A3(g2434C),.A2(g2420C),.A1(g2406C));
AND2_X1 U_g9863C (.ZN(g9863C),.A2(FE_OFN56_g9052C),.A1(g9740C));
AND4_X1 U_I5886C (.ZN(I5886C),.A4(g2254C),.A3(g2249C),.A2(g170C),.A1(g174C));
AND2_X1 U_g6994C (.ZN(g6994C),.A2(FE_OFN141_g3829C),.A1(g6758C));
AND2_X1 U_g9713C (.ZN(g9713C),.A2(FE_OFN63_g9474C),.A1(g1589C));
AND2_X1 U_g4431C (.ZN(g4431C),.A2(g3533C),.A1(g2268C));
AND2_X1 U_g4252C (.ZN(g4252C),.A2(FE_OFN347_g3914C),.A1(g1007C));
AND2_X1 U_g11166C (.ZN(g11166C),.A2(FE_OFN9_g10702C),.A1(g542C));
AND2_X1 U_g7130C (.ZN(g7130C),.A2(g6697C),.A1(g5150C));
AND2_X1 U_g11009C (.ZN(g11009C),.A2(FE_OFN18_g10702C),.A1(g5179C));
AND2_X1 U_g7542C (.ZN(g7542C),.A2(g79C),.A1(FE_OFN85_g2176C));
AND2_X1 U_g8019C (.ZN(g8019C),.A2(FE_OFN310_g4336C),.A1(g6573C));
AND2_X1 U_g11008C (.ZN(g11008C),.A2(FE_OFN18_g10702C),.A1(g5171C));
AND2_X1 U_g3516C (.ZN(g3516C),.A2(FE_OFN298_g3015C),.A1(g1209C));
AND2_X1 U_g8052C (.ZN(g8052C),.A2(FE_OFN305_g5151C),.A1(g7573C));
AND2_X1 U_g3987C (.ZN(g3987C),.A2(FE_OFN359_g18C),.A1(g243C));
AND2_X1 U_g4765C (.ZN(g4765C),.A2(FE_OFN307_g4010C),.A1(g491C));
AND2_X1 U_g11555C (.ZN(g11555C),.A2(FE_OFN27_g11519C),.A1(FE_OFN238_g1781C));
AND2_X1 U_g9857C (.ZN(g9857C),.A2(g9569C),.A1(g9734C));
AND2_X1 U_g8728C (.ZN(g8728C),.A2(g7915C),.A1(g8226C));
AND2_X1 U_g8730C (.ZN(g8730C),.A2(g7917C),.A1(g8230C));
AND2_X1 U_g8185C (.ZN(g8185C),.A2(g8234C),.A1(g664C));
AND2_X1 U_g5194C (.ZN(g5194C),.A2(FE_OFN299_g4457C),.A1(g1610C));
AND2_X1 U_g8385C (.ZN(g8385C),.A2(g8234C),.A1(g5255C));
AND2_X1 U_g4610C (.ZN(g4610C),.A2(g2212C),.A1(g3804C));
AND2_X1 U_g7902C (.ZN(g7902C),.A2(g6449C),.A1(g7661C));
AND2_X1 U_g4073C (.ZN(g4073C),.A2(g3222C),.A1(g3200C));
AND2_X1 U_g8070C (.ZN(g8070C),.A2(FE_OFN198_g7697C),.A1(g682C));
AND2_X1 U_g5731C (.ZN(g5731C),.A2(FE_OFN315_g5117C),.A1(g1583C));
AND2_X1 U_g11238C (.ZN(g11238C),.A2(g11111C),.A1(g4553C));
AND2_X1 U_g4473C (.ZN(g4473C),.A2(FE_OFN302_g3913C),.A1(g1125C));
AND2_X1 U_g8470C (.ZN(g8470C),.A2(FE_OFN210_g7246C),.A1(g8308C));
AND2_X1 U_g5489C (.ZN(g5489C),.A2(FE_OFN358_g3521C),.A1(g557C));
AND2_X1 U_g3991C (.ZN(g3991C),.A2(g2774C),.A1(g1738C));
AND4_X1 U_I5887C (.ZN(I5887C),.A4(g2095C),.A3(g166C),.A2(g2083C),.A1(g2078C));
AND2_X1 U_g7823C (.ZN(g7823C),.A2(FE_OFN209_g6863C),.A1(g1923C));
AND2_X1 U_g4069C (.ZN(g4069C),.A2(g2777C),.A1(g1762C));
AND3_X4 U_g11519C (.ZN(g11519C),.A3(g11492C),.A2(g3015C),.A1(g1317C));
AND2_X1 U_g11176C (.ZN(g11176C),.A2(FE_OFN20_g10702C),.A1(g506C));
AND2_X1 U_g11092C (.ZN(g11092C),.A2(FE_OFN4_g10950C),.A1(g837C));
AND2_X1 U_g11154C (.ZN(g11154C),.A2(FE_OFN278_g10927C),.A1(g330C));
AND2_X1 U_g9608C (.ZN(g9608C),.A2(FE_OFN71_g9292C),.A1(g7C));
AND2_X1 U_g11637C (.ZN(g11637C),.A2(FE_OFN99_g4421C),.A1(g11596C));
AND2_X1 U_g2091C (.ZN(g2091C),.A2(g971C),.A1(g976C));
AND2_X1 U_g8406C (.ZN(g8406C),.A2(g8146C),.A1(g695C));
AND2_X1 U_g5254C (.ZN(g5254C),.A2(FE_OFN357_g3521C),.A1(g549C));
AND2_X1 U_g7260C (.ZN(g7260C),.A2(g2345C),.A1(g6752C));
AND2_X1 U_g5150C (.ZN(g5150C),.A2(g4678C),.A1(g1275C));
AND2_X1 U_g8766C (.ZN(g8766C),.A2(FE_OFN304_g5151C),.A1(g8612C));
AND2_X1 U_g9588C (.ZN(g9588C),.A2(FE_OFN53_g9173C),.A1(g1351C));
AND2_X1 U_g8801C (.ZN(g8801C),.A2(FE_OFN331_g8696C),.A1(g8742C));
AND2_X1 U_g7063C (.ZN(g7063C),.A2(g6586C),.A1(g5008C));
AND2_X1 U_g10303C (.ZN(g10303C),.A2(g9291C),.A1(g9995C));
AND2_X1 U_g5009C (.ZN(g5009C),.A2(FE_OFN154_g4640C),.A1(g1486C));
AND2_X1 U_g9665C (.ZN(g9665C),.A2(FE_OFN48_g9151C),.A1(g1314C));
AND2_X2 U_g8748C (.ZN(g8748C),.A2(g8488C),.A1(I9810C));
AND2_X1 U_g11215C (.ZN(g11215C),.A2(FE_OFN279_g11157C),.A1(g953C));
AND2_X1 U_g10750C (.ZN(g10750C),.A2(FE_OFN102_g3586C),.A1(g10597C));
AND3_X1 U_g5769C (.ZN(g5769C),.A3(g3818C),.A2(FE_OFN200_g4921C),.A1(g3092C));
AND2_X1 U_g6673C (.ZN(g6673C),.A2(I9326C),.A1(g90C));
AND2_X1 U_g5212C (.ZN(g5212C),.A2(g4678C),.A1(g1255C));
AND2_X1 U_g7720C (.ZN(g7720C),.A2(FE_OFN191_g6488C),.A1(g727C));
AND3_X1 U_g5918C (.ZN(g5918C),.A3(g4609C),.A2(FE_OFN184_I7048C),.A1(g109C));
AND2_X1 U_g8045C (.ZN(g8045C),.A2(g5128C),.A1(g7547C));
AND2_X1 U_g8173C (.ZN(g8173C),.A2(FE_OFN363_I5565C),.A1(g7971C));
AND2_X1 U_g11349C (.ZN(g11349C),.A2(g7914C),.A1(g11288C));
AND2_X1 U_g7843C (.ZN(g7843C),.A2(g5919C),.A1(g7599C));
AND2_X1 U_g9696C (.ZN(g9696C),.A2(FE_OFN59_g9432C),.A1(g281C));
AND2_X1 U_g6772C (.ZN(g6772C),.A2(g722C),.A1(g6228C));
AND2_X1 U_g6058C (.ZN(g6058C),.A2(g85C),.A1(g1035C));
AND2_X1 U_g6531C (.ZN(g6531C),.A2(FE_OFN283_I8869C),.A1(g79C));
AND2_X1 U_g6743C (.ZN(g6743C),.A2(FE_OFN219_g5557C),.A1(g4106C));
AND2_X1 U_g6890C (.ZN(g6890C),.A2(g6403C),.A1(g6752C));
AND2_X1 U_g7549C (.ZN(g7549C),.A2(FE_OFN137_g3829C),.A1(g7269C));
AND2_X1 U_g8169C (.ZN(g8169C),.A2(I11360C),.A1(g35C));
AND2_X1 U_g11304C (.ZN(g11304C),.A2(g11243C),.A1(g4585C));
AND2_X1 U_g9944C (.ZN(g9944C),.A2(FE_OFN68_g9392C),.A1(g9924C));
AND2_X4 U_g9240C (.ZN(g9240C),.A2(g8962C),.A1(FE_OFN277_g48C));
AND2_X1 U_g8059C (.ZN(g8059C),.A2(FE_OFN177_g5919C),.A1(g7592C));
AND2_X1 U_g8718C (.ZN(g8718C),.A2(g7903C),.A1(g8203C));
AND2_X1 U_g8767C (.ZN(g8767C),.A2(FE_OFN304_g5151C),.A1(g8616C));
AND2_X1 U_g9316C (.ZN(g9316C),.A2(g48C),.A1(g8877C));
AND2_X1 U_g7625C (.ZN(g7625C),.A2(FE_OFN191_g6488C),.A1(g673C));
AND2_X1 U_g8793C (.ZN(g8793C),.A2(FE_OFN331_g8696C),.A1(g8644C));
AND2_X1 U_g2940C (.ZN(g2940C),.A2(g1654C),.A1(g2424C));
AND2_X1 U_g4114C (.ZN(g4114C),.A2(g3301C),.A1(g1351C));
AND2_X1 U_g11636C (.ZN(g11636C),.A2(g7897C),.A1(g11624C));
AND2_X1 U_g10949C (.ZN(g10949C),.A2(g10809C),.A1(g2947C));
AND2_X1 U_g3563C (.ZN(g3563C),.A2(g2126C),.A1(g3275C));
AND2_X1 U_g10948C (.ZN(g10948C),.A2(g10809C),.A1(g2223C));
AND2_X1 U_g8246C (.ZN(g8246C),.A2(g7438C),.A1(g7846C));
AND2_X1 U_g5788C (.ZN(g5788C),.A2(g5222C),.A1(g1540C));
AND2_X1 U_g4008C (.ZN(g4008C),.A2(FE_OFN224_g2276C),.A1(FE_OFN236_g1776C));
AND2_X1 U_g9596C (.ZN(g9596C),.A2(g9010C),.A1(g928C));
AND2_X1 U_g5249C (.ZN(g5249C),.A2(FE_OFN288_g4263C),.A1(g1089C));
AND2_X1 U_g11585C (.ZN(g11585C),.A2(g11539C),.A1(g1321C));
AND2_X1 U_g3089C (.ZN(g3089C),.A2(g2050C),.A1(g2054C));
AND2_X1 U_g4972C (.ZN(g4972C),.A2(FE_OFN147_g4682C),.A1(g1436C));
AND2_X1 U_g11554C (.ZN(g11554C),.A2(FE_OFN27_g11519C),.A1(g1776C));
AND2_X1 U_g7586C (.ZN(g7586C),.A2(g5420C),.A1(g7096C));
AND2_X1 U_g10673C (.ZN(g10673C),.A2(FE_OFN79_g8700C),.A1(g10417C));
AND3_X1 U_g4806C (.ZN(g4806C),.A3(g2493C),.A2(g3992C),.A1(g3215C));
AND2_X1 U_g5485C (.ZN(g5485C),.A2(FE_OFN333_g4294C),.A1(g1914C));
AND2_X1 U_g9936C (.ZN(g9936C),.A2(FE_OFN60_g9624C),.A1(g9915C));
AND2_X1 U_g2910C (.ZN(g2910C),.A2(g1660C),.A1(g2424C));
AND2_X1 U_g9317C (.ZN(g9317C),.A2(g8875C),.A1(g6109C));
AND2_X1 U_g10933C (.ZN(g10933C),.A2(g3982C),.A1(g10853C));
AND2_X1 U_g8388C (.ZN(g8388C),.A2(g7246C),.A1(g8177C));
AND2_X1 U_g4465C (.ZN(g4465C),.A2(FE_OFN302_g3913C),.A1(g1117C));
AND2_X1 U_g7141C (.ZN(g7141C),.A2(g6716C),.A1(g5230C));
AND2_X1 U_g10508C (.ZN(g10508C),.A2(FE_OFN336_g1690C),.A1(g10013C));
AND2_X1 U_g4230C (.ZN(g4230C),.A2(FE_OFN132_g3015C),.A1(g1095C));
AND2_X1 U_g10634C (.ZN(g10634C),.A2(g3829C),.A1(g10382C));
AND2_X1 U_g9601C (.ZN(g9601C),.A2(g9192C),.A1(g922C));
AND2_X1 U_g6126C (.ZN(g6126C),.A2(FE_OFN322_g4449C),.A1(g3681C));
AND2_X1 U_g6326C (.ZN(g6326C),.A2(FE_OFN115_g4807C),.A1(g1250C));
AND2_X1 U_g7710C (.ZN(g7710C),.A2(FE_OFN191_g6488C),.A1(g700C));
AND2_X1 U_g8028C (.ZN(g8028C),.A2(g7438C),.A1(g7375C));
AND2_X1 U_g6760C (.ZN(g6760C),.A2(g6221C),.A1(g786C));
AND2_X1 U_g5640C (.ZN(g5640C),.A2(FE_OFN290_g4880C),.A1(g1059C));
AND2_X1 U_g5031C (.ZN(g5031C),.A2(FE_OFN153_g4640C),.A1(g1478C));
AND2_X1 U_g4550C (.ZN(g4550C),.A2(FE_OFN344_g3586C),.A1(g342C));
AND2_X1 U_g7879C (.ZN(g7879C),.A2(FE_OFN366_g3521C),.A1(g5286C));
AND2_X1 U_g7962C (.ZN(g7962C),.A2(g6403C),.A1(g7730C));
AND2_X1 U_g9597C (.ZN(g9597C),.A2(FE_OFN46_g9125C),.A1(g1170C));
AND2_X1 U_g10452C (.ZN(g10452C),.A2(FE_OFN234_g2024C),.A1(g10439C));
AND2_X1 U_g4891C (.ZN(g4891C),.A2(g4739C),.A1(g631C));
AND2_X1 U_g5005C (.ZN(g5005C),.A2(FE_OFN154_g4640C),.A1(g1490C));
AND2_X1 U_g6423C (.ZN(g6423C),.A2(FE_OFN217_g5013C),.A1(g4348C));
AND2_X1 U_g8108C (.ZN(g8108C),.A2(g7952C),.A1(g1891C));
AND3_X4 U_g4807C (.ZN(g4807C),.A3(I6360C),.A2(g1289C),.A1(g3015C));
AND2_X1 U_g5911C (.ZN(g5911C),.A2(g4977C),.A1(g3322C));
AND2_X1 U_g9937C (.ZN(g9937C),.A2(FE_OFN60_g9624C),.A1(g9916C));
AND2_X1 U_g9840C (.ZN(g9840C),.A2(g9747C),.A1(g9704C));
AND2_X1 U_g10780C (.ZN(g10780C),.A2(g4467C),.A1(g10723C));
AND2_X1 U_g8217C (.ZN(g8217C),.A2(g7883C),.A1(g1872C));
AND2_X1 U_g11013C (.ZN(g11013C),.A2(FE_OFN18_g10702C),.A1(g5209C));
AND2_X1 U_g9390C (.ZN(g9390C),.A2(FE_OFN48_g9151C),.A1(g1333C));
AND2_X1 U_g11214C (.ZN(g11214C),.A2(FE_OFN279_g11157C),.A1(g950C));
AND2_X1 U_g6327C (.ZN(g6327C),.A2(FE_OFN115_g4807C),.A1(g1255C));
AND2_X1 U_g4342C (.ZN(g4342C),.A2(FE_OFN351_g3913C),.A1(g1149C));
AND2_X1 U_g5796C (.ZN(g5796C),.A2(FE_OFN321_g5261C),.A1(g1564C));
AND2_X1 U_g5473C (.ZN(g5473C),.A2(FE_OFN367_g3521C),.A1(g546C));
AND2_X1 U_g6346C (.ZN(g6346C),.A2(g5878C),.A1(g5038C));
AND2_X1 U_g6633C (.ZN(g6633C),.A2(FE_OFN282_g6165C),.A1(g354C));
AND2_X1 U_g11005C (.ZN(g11005C),.A2(FE_OFN13_g10702C),.A1(g5119C));
AND2_X1 U_g8365C (.ZN(g8365C),.A2(g8146C),.A1(g668C));
AND2_X1 U_g8048C (.ZN(g8048C),.A2(g5919C),.A1(g7558C));
AND2_X1 U_g4481C (.ZN(g4481C),.A2(g3906C),.A1(g1713C));
AND2_X1 U_g4097C (.ZN(g4097C),.A2(g3060C),.A1(g2677C));
AND2_X1 U_g8055C (.ZN(g8055C),.A2(FE_OFN305_g5151C),.A1(g7588C));
AND2_X1 U_g4497C (.ZN(g4497C),.A2(FE_OFN344_g3586C),.A1(g351C));
AND2_X1 U_g9942C (.ZN(g9942C),.A2(FE_OFN67_g9367C),.A1(g9922C));
AND2_X1 U_g6696C (.ZN(g6696C),.A2(I9326C),.A1(g94C));
AND3_X1 U_g10731C (.ZN(g10731C),.A3(g10665C),.A2(g1850C),.A1(g5118C));
AND2_X1 U_g8827C (.ZN(g8827C),.A2(g8696C),.A1(g8552C));
AND2_X1 U_g5540C (.ZN(g5540C),.A2(g4292C),.A1(g1727C));
AND2_X1 U_g4960C (.ZN(g4960C),.A2(FE_OFN147_g4682C),.A1(g1403C));
AND2_X1 U_g8846C (.ZN(g8846C),.A2(FE_OFN328_g8709C),.A1(g8615C));
AND2_X1 U_g6508C (.ZN(g6508C),.A2(FE_OFN363_I5565C),.A1(g5983C));
AND2_X1 U_g6240C (.ZN(g6240C),.A2(g5361C),.A1(g182C));
AND2_X1 U_g7931C (.ZN(g7931C),.A2(g7446C),.A1(g52C));
AND2_X1 U_g5287C (.ZN(g5287C),.A2(g4782C),.A1(I6260C));
AND2_X1 U_g6472C (.ZN(g6472C),.A2(g1936C),.A1(g5853C));
AND2_X1 U_g11100C (.ZN(g11100C),.A2(FE_OFN4_g10950C),.A1(g853C));
AND2_X1 U_g11235C (.ZN(g11235C),.A2(g11107C),.A1(g4529C));
AND2_X1 U_g5199C (.ZN(g5199C),.A2(FE_OFN288_g4263C),.A1(g1068C));
AND2_X1 U_g6316C (.ZN(g6316C),.A2(FE_OFN117_g4807C),.A1(g1270C));
AND2_X1 U_g7515C (.ZN(g7515C),.A2(g70C),.A1(FE_OFN85_g2176C));
AND2_X1 U_g10583C (.ZN(g10583C),.A2(g10515C),.A1(g10518C));
AND2_X1 U_g5781C (.ZN(g5781C),.A2(g5222C),.A1(g1537C));
AND2_X1 U_g8018C (.ZN(g8018C),.A2(g7438C),.A1(g7742C));
AND2_X1 U_g4401C (.ZN(g4401C),.A2(g3772C),.A1(g1845C));
AND3_X1 U_g8994C (.ZN(g8994C),.A3(g8783C),.A2(FE_OFN92_g2216C),.A1(g8110C));
AND2_X1 U_g2950C (.ZN(g2950C),.A2(g1666C),.A1(g2424C));
AND2_X1 U_g5510C (.ZN(g5510C),.A2(g4289C),.A1(g1630C));
AND2_X1 U_g6347C (.ZN(g6347C),.A2(FE_OFN320_g5361C),.A1(g275C));
AND2_X1 U_g9357C (.ZN(g9357C),.A2(g9223C),.A1(g962C));
AND2_X1 U_g4828C (.ZN(g4828C),.A2(g695C),.A1(g4106C));
AND2_X1 U_g11407C (.ZN(g11407C),.A2(g4807C),.A1(g11249C));
AND2_X1 U_g4727C (.ZN(g4727C),.A2(FE_OFN300_g4002C),.A1(g386C));
AND2_X1 U_g10357C (.ZN(g10357C),.A2(FE_OFN269_g109C),.A1(I15500C));
AND2_X1 U_g10743C (.ZN(g10743C),.A2(FE_OFN364_g3015C),.A1(g10639C));
AND2_X1 U_g5259C (.ZN(g5259C),.A2(g4739C),.A1(g627C));
AND2_X1 U_g5694C (.ZN(g5694C),.A2(FE_OFN365_g5361C),.A1(g162C));
AND2_X1 U_g10769C (.ZN(g10769C),.A2(FE_OFN297_g3015C),.A1(g10652C));
AND2_X1 U_g11584C (.ZN(g11584C),.A2(g11539C),.A1(g1318C));
AND2_X1 U_g4932C (.ZN(g4932C),.A2(FE_OFN290_g4880C),.A1(g1065C));
AND2_X1 U_g10768C (.ZN(g10768C),.A2(FE_OFN293_g3015C),.A1(g10649C));
AND2_X1 U_g6820C (.ZN(g6820C),.A2(FE_OFN178_g5354C),.A1(g1362C));
AND2_X1 U_g4068C (.ZN(g4068C),.A2(FE_OFN224_g2276C),.A1(FE_OFN251_g1801C));
AND2_X1 U_g6317C (.ZN(g6317C),.A2(FE_OFN117_g4807C),.A1(g1304C));
AND2_X1 U_g5215C (.ZN(g5215C),.A2(g3275C),.A1(g4276C));
AND2_X1 U_g4576C (.ZN(g4576C),.A2(g4010C),.A1(g530C));
AND2_X1 U_g6775C (.ZN(g6775C),.A2(g6231C),.A1(g822C));
AND2_X4 U_g3829C (.ZN(g3829C),.A2(g1696C),.A1(g2028C));
AND2_X1 U_g10662C (.ZN(g10662C),.A2(g10396C),.A1(g8700C));
AND2_X1 U_g8101C (.ZN(g8101C),.A2(FE_OFN207_g6863C),.A1(g5484C));
AND2_X1 U_g5825C (.ZN(g5825C),.A2(g5318C),.A1(g3204C));
AND4_X1 U_I6310C (.ZN(I6310C),.A4(g2435C),.A3(g2421C),.A2(g2407C),.A1(g2396C));
AND2_X1 U_g7884C (.ZN(g7884C),.A2(FE_OFN334_g7045C),.A1(g7457C));
AND2_X1 U_g5008C (.ZN(g5008C),.A2(FE_OFN303_g4678C),.A1(g1292C));
AND2_X1 U_g3974C (.ZN(g3974C),.A2(FE_OFN260_g18C),.A1(g231C));
AND2_X1 U_g9949C (.ZN(g9949C),.A2(FE_OFN68_g9392C),.A1(g9929C));
AND2_X1 U_g2531C (.ZN(g2531C),.A2(g668C),.A1(g658C));
AND2_X2 U_g9292C (.ZN(g9292C),.A2(g48C),.A1(g8878C));
AND2_X1 U_g10778C (.ZN(g10778C),.A2(g10679C),.A1(g1027C));
AND2_X1 U_g8041C (.ZN(g8041C),.A2(g5128C),.A1(g7524C));
AND2_X1 U_g6079C (.ZN(g6079C),.A2(FE_OFN273_g85C),.A1(g1053C));
AND2_X1 U_g7235C (.ZN(g7235C),.A2(g6447C),.A1(g6663C));
AND2_X1 U_g9603C (.ZN(g9603C),.A2(FE_OFN46_g9125C),.A1(g1173C));
AND2_X1 U_g6840C (.ZN(g6840C),.A2(FE_OFN180_g5354C),.A1(g248C));
AND2_X1 U_g9850C (.ZN(g9850C),.A2(g9579C),.A1(g9726C));
AND2_X1 U_g7988C (.ZN(g7988C),.A2(g7379C),.A1(g1878C));
AND2_X1 U_g5228C (.ZN(g5228C),.A2(FE_OFN288_g4263C),.A1(g1086C));
AND2_X1 U_g7134C (.ZN(g7134C),.A2(g6354C),.A1(g5587C));
AND2_X1 U_g5934C (.ZN(g5934C),.A2(g1965C),.A1(g5215C));
AND2_X1 U_g5230C (.ZN(g5230C),.A2(g4678C),.A1(g1265C));
AND2_X1 U_g8168C (.ZN(g8168C),.A2(FE_OFN89_I11360C),.A1(g34C));
AND2_X1 U_g9583C (.ZN(g9583C),.A2(g8995C),.A1(g886C));
AND2_X1 U_g10672C (.ZN(g10672C),.A2(g9473C),.A1(g10414C));
AND2_X1 U_g3287C (.ZN(g3287C),.A2(g5188C),.A1(g802C));
AND2_X1 U_g8772C (.ZN(g8772C),.A2(FE_OFN304_g5151C),.A1(g8627C));
AND2_X1 U_g4893C (.ZN(g4893C),.A2(g4739C),.A1(g635C));
AND2_X1 U_g10331C (.ZN(g10331C),.A2(FE_OFN269_g109C),.A1(I15510C));
AND2_X1 U_g8505C (.ZN(g8505C),.A2(FE_OFN359_g18C),.A1(g8309C));
AND2_X1 U_g10449C (.ZN(g10449C),.A2(FE_OFN235_g2024C),.A1(g10433C));
AND2_X1 U_g11273C (.ZN(g11273C),.A2(g11199C),.A1(g4765C));
AND2_X1 U_g8734C (.ZN(g8734C),.A2(g7923C),.A1(g8187C));
AND2_X1 U_g5913C (.ZN(g5913C),.A2(g85C),.A1(g1041C));
AND2_X1 U_g10448C (.ZN(g10448C),.A2(FE_OFN235_g2024C),.A1(g10421C));
AND2_X1 U_g6163C (.ZN(g6163C),.A2(g5354C),.A1(g4572C));
AND2_X1 U_g6363C (.ZN(g6363C),.A2(FE_OFN320_g5361C),.A1(g284C));
AND2_X1 U_g7202C (.ZN(g7202C),.A2(FE_OFN322_g4449C),.A1(g5226C));
AND2_X1 U_g11463C (.ZN(g11463C),.A2(FE_OFN99_g4421C),.A1(g11229C));
AND2_X1 U_g8074C (.ZN(g8074C),.A2(FE_OFN198_g7697C),.A1(g718C));
AND2_X1 U_g4325C (.ZN(g4325C),.A2(FE_OFN351_g3913C),.A1(g1166C));
AND2_X1 U_g8474C (.ZN(g8474C),.A2(g5521C),.A1(g8383C));
AND2_X1 U_g11234C (.ZN(g11234C),.A2(g11107C),.A1(g4518C));
AND2_X1 U_g5266C (.ZN(g5266C),.A2(FE_OFN335_g4737C),.A1(g718C));
AND2_X1 U_g4483C (.ZN(g4483C),.A2(FE_OFN103_g3586C),.A1(g336C));
AND2_X1 U_g5248C (.ZN(g5248C),.A2(FE_OFN335_g4737C),.A1(g673C));
AND2_X1 U_g11514C (.ZN(g11514C),.A2(FE_OFN176_g5151C),.A1(g11491C));
AND2_X1 U_g5255C (.ZN(g5255C),.A2(FE_OFN335_g4737C),.A1(g682C));
AND2_X1 U_g4106C (.ZN(g4106C),.A2(g686C),.A1(g3284C));
AND2_X1 U_g2760C (.ZN(g2760C),.A2(g2091C),.A1(g981C));
AND2_X1 U_g5097C (.ZN(g5097C),.A2(g4608C),.A1(g1786C));
AND2_X1 U_g5726C (.ZN(g5726C),.A2(FE_OFN315_g5117C),.A1(g1601C));
AND2_X1 U_g5497C (.ZN(g5497C),.A2(FE_OFN357_g3521C),.A1(g560C));
AND2_X4 U_g5354C (.ZN(g5354C),.A2(I7048C),.A1(FE_OFN352_g109C));
AND2_X1 U_g7933C (.ZN(g7933C),.A2(g7450C),.A1(g55C));
AND2_X1 U_g9617C (.ZN(g9617C),.A2(g9274C),.A1(g9C));
AND2_X1 U_g9906C (.ZN(g9906C),.A2(g9680C),.A1(g9873C));
AND2_X1 U_g11012C (.ZN(g11012C),.A2(FE_OFN18_g10702C),.A1(g5196C));
AND2_X1 U_g7050C (.ZN(g7050C),.A2(g6702C),.A1(g5001C));
AND2_X1 U_g10971C (.ZN(g10971C),.A2(g2045C),.A1(g10849C));
AND2_X1 U_g4904C (.ZN(g4904C),.A2(g4243C),.A1(g1850C));
AND2_X1 U_g10369C (.ZN(g10369C),.A2(FE_OFN235_g2024C),.A1(g10361C));
AND2_X1 U_g8400C (.ZN(g8400C),.A2(g8234C),.A1(g5271C));
AND2_X1 U_g4345C (.ZN(g4345C),.A2(FE_OFN289_g4679C),.A1(g1169C));
AND2_X1 U_g2161C (.ZN(g2161C),.A2(I5085C),.A1(I5084C));
AND2_X1 U_g5001C (.ZN(g5001C),.A2(FE_OFN303_g4678C),.A1(g1300C));
AND2_X1 U_g9945C (.ZN(g9945C),.A2(FE_OFN68_g9392C),.A1(g9925C));
AND2_X1 U_g7271C (.ZN(g7271C),.A2(g6354C),.A1(g5028C));
AND2_X1 U_g9709C (.ZN(g9709C),.A2(FE_OFN70_g9490C),.A1(g1524C));
AND2_X1 U_g4223C (.ZN(g4223C),.A2(FE_OFN347_g3914C),.A1(g1003C));
AND2_X1 U_g10716C (.ZN(g10716C),.A2(g10396C),.A1(g10497C));
AND2_X1 U_g11291C (.ZN(g11291C),.A2(g4379C),.A1(g11247C));
AND2_X1 U_g6661C (.ZN(g6661C),.A2(FE_OFN97_I8869C),.A1(g73C));
AND2_X1 U_g11173C (.ZN(g11173C),.A2(FE_OFN21_g10702C),.A1(g491C));
AND2_X1 U_g6075C (.ZN(g6075C),.A2(g5613C),.A1(g549C));
AND2_X1 U_g8023C (.ZN(g8023C),.A2(g7438C),.A1(g7367C));
AND2_X1 U_g9907C (.ZN(g9907C),.A2(g9680C),.A1(g9888C));
AND2_X1 U_g10582C (.ZN(g10582C),.A2(g9473C),.A1(g10339C));
AND2_X1 U_g5746C (.ZN(g5746C),.A2(FE_OFN353_g5117C),.A1(g1589C));
AND2_X1 U_g5221C (.ZN(g5221C),.A2(g4678C),.A1(g1260C));
AND2_X1 U_g9959C (.ZN(g9959C),.A2(FE_OFN280_g9536C),.A1(g9950C));
AND2_X1 U_g7674C (.ZN(g7674C),.A2(g3880C),.A1(g5857C));
AND2_X1 U_g9690C (.ZN(g9690C),.A2(g9432C),.A1(g266C));
AND2_X1 U_g6627C (.ZN(g6627C),.A2(FE_OFN283_I8869C),.A1(g58C));
AND2_X1 U_g5703C (.ZN(g5703C),.A2(FE_OFN365_g5361C),.A1(g174C));
AND2_X1 U_g4522C (.ZN(g4522C),.A2(FE_OFN344_g3586C),.A1(g360C));
AND2_X1 U_g4115C (.ZN(g4115C),.A2(g3060C),.A1(FE_OFN236_g1776C));
AND2_X1 U_g7541C (.ZN(g7541C),.A2(I6360C),.A1(g7075C));
AND2_X1 U_g10627C (.ZN(g10627C),.A2(FE_OFN227_g3880C),.A1(g10452C));
AND2_X1 U_g4047C (.ZN(g4047C),.A2(FE_OFN225_g2276C),.A1(FE_OFN238_g1781C));
AND2_X1 U_g6526C (.ZN(g6526C),.A2(FE_OFN283_I8869C),.A1(g76C));
AND2_X1 U_g2944C (.ZN(g2944C),.A2(g1669C),.A1(g2424C));
AND2_X1 U_g6646C (.ZN(g6646C),.A2(g6165C),.A1(g360C));
AND2_X1 U_g7132C (.ZN(g7132C),.A2(g6702C),.A1(g5182C));
AND2_X1 U_g11029C (.ZN(g11029C),.A2(FE_OFN17_g10702C),.A1(g401C));
AND2_X1 U_g8051C (.ZN(g8051C),.A2(FE_OFN305_g5151C),.A1(g7572C));
AND2_X1 U_g8127C (.ZN(g8127C),.A2(g7949C),.A1(g1927C));
AND2_X1 U_g7209C (.ZN(g7209C),.A2(g6432C),.A1(g3804C));
AND2_X1 U_g11028C (.ZN(g11028C),.A2(FE_OFN17_g10702C),.A1(g396C));
AND2_X1 U_g6439C (.ZN(g6439C),.A2(g5919C),.A1(g3631C));
AND2_X1 U_g10742C (.ZN(g10742C),.A2(g3586C),.A1(g10655C));
AND2_X1 U_g9110C (.ZN(g9110C),.A2(FE_OFN359_g18C),.A1(g8880C));
AND2_X1 U_g10681C (.ZN(g10681C),.A2(g3586C),.A1(g10567C));
AND2_X1 U_g4537C (.ZN(g4537C),.A2(g4002C),.A1(g444C));
AND2_X1 U_g9663C (.ZN(g9663C),.A2(FE_OFN39_g9223C),.A1(g959C));
AND2_X1 U_g5349C (.ZN(g5349C),.A2(g4617C),.A1(g2126C));
AND2_X1 U_g8732C (.ZN(g8732C),.A2(g7919C),.A1(g8200C));
AND2_X1 U_g3807C (.ZN(g3807C),.A2(g3062C),.A1(g3003C));
AND2_X1 U_g5848C (.ZN(g5848C),.A2(g5519C),.A1(g3860C));
AND2_X1 U_g8508C (.ZN(g8508C),.A2(FE_OFN330_g7638C),.A1(g8411C));
AND2_X1 U_g8072C (.ZN(g8072C),.A2(FE_OFN199_g7697C),.A1(g700C));
AND2_X1 U_g5699C (.ZN(g5699C),.A2(g5117C),.A1(g1592C));
AND2_X1 U_g11240C (.ZN(g11240C),.A2(g11111C),.A1(g4560C));
AND2_X1 U_g5398C (.ZN(g5398C),.A2(g2224C),.A1(g4610C));
AND2_X1 U_g6616C (.ZN(g6616C),.A2(FE_OFN363_I5565C),.A1(g6105C));
AND2_X1 U_g10690C (.ZN(g10690C),.A2(FE_OFN136_g3863C),.A1(g10387C));
AND2_X1 U_g8043C (.ZN(g8043C),.A2(FE_OFN305_g5151C),.A1(g7582C));
AND2_X1 U_g9590C (.ZN(g9590C),.A2(g8995C),.A1(g895C));
AND2_X1 U_g4128C (.ZN(g4128C),.A2(g627C),.A1(g1976C));
AND2_X1 U_g6404C (.ZN(g6404C),.A2(FE_OFN217_g5013C),.A1(g2132C));
AND2_X1 U_g6647C (.ZN(g6647C),.A2(g5808C),.A1(g87C));
AND2_X1 U_g10504C (.ZN(g10504C),.A2(FE_OFN336_g1690C),.A1(g10001C));
AND2_X1 U_g9657C (.ZN(g9657C),.A2(g9205C),.A1(g919C));
AND2_X1 U_g4542C (.ZN(g4542C),.A2(FE_OFN344_g3586C),.A1(g366C));
AND2_X1 U_g4330C (.ZN(g4330C),.A2(FE_OFN351_g3913C),.A1(g1163C));
AND2_X1 U_g3497C (.ZN(g3497C),.A2(g1900C),.A1(g2804C));
AND2_X1 U_g5524C (.ZN(g5524C),.A2(g3906C),.A1(g1678C));
AND2_X1 U_g8147C (.ZN(g8147C),.A2(g7907C),.A1(g928C));
AND2_X1 U_g4554C (.ZN(g4554C),.A2(g4010C),.A1(g542C));
AND2_X1 U_g9899C (.ZN(g9899C),.A2(g9367C),.A1(g9713C));
AND2_X1 U_g5258C (.ZN(g5258C),.A2(FE_OFN335_g4737C),.A1(g700C));
AND2_X1 U_g7736C (.ZN(g7736C),.A2(FE_OFN226_g3880C),.A1(g5814C));
AND2_X1 U_g6224C (.ZN(g6224C),.A2(FE_OFN306_g5128C),.A1(g1520C));
AND2_X1 U_g10626C (.ZN(g10626C),.A2(FE_OFN369_g4525C),.A1(g10453C));
AND2_X1 U_g6320C (.ZN(g6320C),.A2(FE_OFN118_g4807C),.A1(g1292C));
AND2_X1 U_g7623C (.ZN(g7623C),.A2(FE_OFN191_g6488C),.A1(g664C));
AND2_X1 U_g10299C (.ZN(g10299C),.A2(g10013C),.A1(FE_OFN76_g8700C));
AND2_X1 U_g7889C (.ZN(g7889C),.A2(g3814C),.A1(g5304C));
AND2_X1 U_g10298C (.ZN(g10298C),.A2(g10007C),.A1(g8700C));
AND2_X1 U_g8413C (.ZN(g8413C),.A2(g8146C),.A1(g722C));
AND2_X1 U_g3979C (.ZN(g3979C),.A2(FE_OFN260_g18C),.A1(g237C));
AND2_X1 U_g4902C (.ZN(g4902C),.A2(g4243C),.A1(g1848C));
AND2_X1 U_g5211C (.ZN(g5211C),.A2(FE_OFN288_g4263C),.A1(g1080C));
AND2_X1 U_g4512C (.ZN(g4512C),.A2(FE_OFN344_g3586C),.A1(g357C));
AND2_X1 U_g7722C (.ZN(g7722C),.A2(g6449C),.A1(g7127C));
AND2_X1 U_g9844C (.ZN(g9844C),.A2(g9522C),.A1(g9714C));
AND2_X1 U_g4490C (.ZN(g4490C),.A2(FE_OFN302_g3913C),.A1(g1141C));
AND2_X1 U_g6516C (.ZN(g6516C),.A2(FE_OFN363_I5565C),.A1(g5993C));
AND2_X1 U_g5026C (.ZN(g5026C),.A2(FE_OFN153_g4640C),.A1(g1453C));
AND2_X1 U_g8820C (.ZN(g8820C),.A2(g4737C),.A1(g8705C));
AND2_X1 U_g10737C (.ZN(g10737C),.A2(FE_OFN133_g3015C),.A1(g10597C));
AND3_X1 U_g8936C (.ZN(g8936C),.A3(g8849C),.A2(FE_OFN93_g2216C),.A1(g8115C));
AND2_X1 U_g10232C (.ZN(g10232C),.A2(g9974C),.A1(FE_OFN76_g8700C));
AND2_X1 U_g6771C (.ZN(g6771C),.A2(FE_OFN320_g5361C),.A1(g263C));
AND2_X1 U_g5170C (.ZN(g5170C),.A2(g4457C),.A1(g1811C));
AND2_X1 U_g8117C (.ZN(g8117C),.A2(FE_OFN207_g6863C),.A1(g5514C));
AND2_X1 U_g4529C (.ZN(g4529C),.A2(g4002C),.A1(g448C));
AND2_X1 U_g4348C (.ZN(g4348C),.A2(g1909C),.A1(g3497C));
AND2_X1 U_g9966C (.ZN(g9966C),.A2(FE_OFN280_g9536C),.A1(g9956C));
AND2_X1 U_g5280C (.ZN(g5280C),.A2(g2118C),.A1(g3967C));
AND2_X1 U_g7139C (.ZN(g7139C),.A2(g6716C),.A1(g5212C));
AND2_X1 U_g11099C (.ZN(g11099C),.A2(g10883C),.A1(g382C));
AND2_X1 U_g6892C (.ZN(g6892C),.A2(g5013C),.A1(g6472C));
AND2_X1 U_g9705C (.ZN(g9705C),.A2(g9474C),.A1(g1580C));
AND2_X1 U_g10512C (.ZN(g10512C),.A2(FE_OFN336_g1690C),.A1(g10025C));
AND2_X1 U_g11098C (.ZN(g11098C),.A2(FE_OFN4_g10950C),.A1(g849C));
AND2_X1 U_g8775C (.ZN(g8775C),.A2(FE_OFN304_g5151C),.A1(g8628C));
AND2_X1 U_g5083C (.ZN(g5083C),.A2(g4782C),.A1(g2510C));
AND2_X1 U_g5544C (.ZN(g5544C),.A2(FE_OFN291_g4880C),.A1(g1687C));
AND2_X1 U_g11272C (.ZN(g11272C),.A2(g11199C),.A1(g4760C));
AND2_X1 U_g5483C (.ZN(g5483C),.A2(g3906C),.A1(g1621C));
AND2_X1 U_g9948C (.ZN(g9948C),.A2(FE_OFN68_g9392C),.A1(g9928C));
AND2_X1 U_g4063C (.ZN(g4063C),.A2(FE_OFN224_g2276C),.A1(FE_OFN239_g1796C));
AND2_X1 U_g11462C (.ZN(g11462C),.A2(FE_OFN99_g4421C),.A1(g11227C));
AND2_X1 U_g6738C (.ZN(g6738C),.A2(FE_OFN219_g5557C),.A1(g2531C));
AND2_X1 U_g8060C (.ZN(g8060C),.A2(FE_OFN177_g5919C),.A1(g7593C));
AND2_X1 U_g6244C (.ZN(g6244C),.A2(FE_OFN306_g5128C),.A1(g1411C));
AND2_X1 U_g11032C (.ZN(g11032C),.A2(FE_OFN14_g10702C),.A1(g416C));
AND2_X1 U_g10445C (.ZN(g10445C),.A2(g1690C),.A1(g9974C));
AND2_X1 U_g9150C (.ZN(g9150C),.A2(FE_OFN325_g18C),.A1(g8882C));
AND2_X1 U_g10316C (.ZN(g10316C),.A2(g9097C),.A1(g10025C));
AND2_X1 U_g5756C (.ZN(g5756C),.A2(g5261C),.A1(g1531C));
AND2_X1 U_g4720C (.ZN(g4720C),.A2(g4673C),.A1(g1023C));
AND2_X1 U_g9409C (.ZN(g9409C),.A2(g9052C),.A1(g1721C));
AND2_X4 U_g8995C (.ZN(g8995C),.A2(g8929C),.A1(FE_OFN277_g48C));
AND2_X1 U_g6876C (.ZN(g6876C),.A2(g6557C),.A1(g4070C));
AND2_X1 U_g4989C (.ZN(g4989C),.A2(FE_OFN146_g4682C),.A1(g1424C));
AND2_X1 U_g9836C (.ZN(g9836C),.A2(FE_OFN34_g9785C),.A1(g9737C));
AND3_X1 U_g6656C (.ZN(g6656C),.A3(FE_OFN184_I7048C),.A2(g6061C),.A1(g109C));
AND2_X1 U_g5514C (.ZN(g5514C),.A2(FE_OFN333_g4294C),.A1(g1941C));
AND2_X1 U_g8390C (.ZN(g8390C),.A2(g6465C),.A1(g8268C));
AND2_X1 U_g5003C (.ZN(g5003C),.A2(FE_OFN154_g4640C),.A1(g1466C));
AND2_X1 U_g9967C (.ZN(g9967C),.A2(FE_OFN280_g9536C),.A1(g9957C));
AND2_X1 U_g5145C (.ZN(g5145C),.A2(g4673C),.A1(g1639C));
AND2_X1 U_g4971C (.ZN(g4971C),.A2(FE_OFN146_g4682C),.A1(g1419C));
AND2_X1 U_g10753C (.ZN(g10753C),.A2(FE_OFN133_g3015C),.A1(g10649C));
AND2_X1 U_g5695C (.ZN(g5695C),.A2(FE_OFN356_g5361C),.A1(g166C));
AND2_X1 U_g7613C (.ZN(g7613C),.A2(g5013C),.A1(g6940C));
AND2_X1 U_g10736C (.ZN(g10736C),.A2(FE_OFN293_g3015C),.A1(g10658C));
AND2_X1 U_g11220C (.ZN(g11220C),.A2(FE_OFN279_g11157C),.A1(g962C));
AND2_X1 U_g7444C (.ZN(g7444C),.A2(g5557C),.A1(g7277C));
AND2_X1 U_g5536C (.ZN(g5536C),.A2(FE_OFN310_g4336C),.A1(g2970C));
AND2_X1 U_g6663C (.ZN(g6663C),.A2(g2237C),.A1(g6064C));
AND2_X1 U_g4670C (.ZN(g4670C),.A2(g2355C),.A1(g192C));
AND2_X1 U_g6824C (.ZN(g6824C),.A2(FE_OFN178_g5354C),.A1(g1371C));
AND2_X1 U_g4253C (.ZN(g4253C),.A2(FE_OFN132_g3015C),.A1(g1074C));
AND2_X1 U_g8250C (.ZN(g8250C),.A2(g7907C),.A1(g932C));
AND2_X1 U_g8163C (.ZN(g8163C),.A2(g3737C),.A1(g7960C));
AND2_X1 U_g10764C (.ZN(g10764C),.A2(FE_OFN345_g3015C),.A1(g10643C));
AND2_X1 U_g5757C (.ZN(g5757C),.A2(g5222C),.A1(g1552C));
AND2_X1 U_g8032C (.ZN(g8032C),.A2(g7438C),.A1(g7385C));
AND2_X1 U_g11591C (.ZN(g11591C),.A2(g11561C),.A1(g2988C));
AND2_X1 U_g8053C (.ZN(g8053C),.A2(FE_OFN177_g5919C),.A1(g7583C));
AND2_X1 U_g11147C (.ZN(g11147C),.A2(FE_OFN278_g10927C),.A1(g321C));
AND2_X1 U_g5522C (.ZN(g5522C),.A2(g4289C),.A1(g1633C));
AND2_X1 U_g5115C (.ZN(g5115C),.A2(g4572C),.A1(g1394C));
AND2_X1 U_g9837C (.ZN(g9837C),.A2(g9751C),.A1(g9697C));
AND2_X1 U_g9620C (.ZN(g9620C),.A2(FE_OFN40_g9240C),.A1(g976C));
AND2_X1 U_g11151C (.ZN(g11151C),.A2(FE_OFN278_g10927C),.A1(g327C));
AND2_X1 U_g11172C (.ZN(g11172C),.A2(FE_OFN21_g10702C),.A1(g486C));
AND2_X1 U_g7885C (.ZN(g7885C),.A2(g3814C),.A1(g5300C));
AND2_X1 U_g6064C (.ZN(g6064C),.A2(g2230C),.A1(g5398C));
AND3_X1 U_g8929C (.ZN(g8929C),.A3(g8828C),.A2(FE_OFN95_g2216C),.A1(g8095C));
AND2_X1 U_g5595C (.ZN(g5595C),.A2(FE_OFN367_g3521C),.A1(g1621C));
AND2_X1 U_g5537C (.ZN(g5537C),.A2(g4449C),.A1(g2260C));
AND2_X1 U_g9842C (.ZN(g9842C),.A2(g9516C),.A1(g9708C));
AND2_X1 U_g4141C (.ZN(g4141C),.A2(g3060C),.A1(FE_OFN252_g1791C));
AND2_X1 U_g4341C (.ZN(g4341C),.A2(FE_OFN103_g3586C),.A1(g339C));
AND2_X4 U_g9192C (.ZN(g9192C),.A2(g8955C),.A1(FE_OFN277_g48C));
AND2_X1 U_g7679C (.ZN(g7679C),.A2(g6863C),.A1(g1950C));
AND2_X1 U_g7378C (.ZN(g7378C),.A2(FE_OFN226_g3880C),.A1(g5847C));
AND2_X1 U_g5612C (.ZN(g5612C),.A2(FE_OFN357_g3521C),.A1(g1627C));
AND2_X1 U_g7135C (.ZN(g7135C),.A2(g6355C),.A1(g869C));
AND2_X1 U_g10970C (.ZN(g10970C),.A2(g3390C),.A1(g10852C));
AND2_X1 U_g11025C (.ZN(g11025C),.A2(FE_OFN9_g10702C),.A1(g426C));
AND2_X1 U_g9854C (.ZN(g9854C),.A2(g9563C),.A1(g9730C));
AND2_X1 U_g7182C (.ZN(g7182C),.A2(FE_OFN213_g6003C),.A1(g1878C));
AND2_X1 U_g9941C (.ZN(g9941C),.A2(FE_OFN67_g9367C),.A1(g9921C));
AND2_X1 U_g6194C (.ZN(g6194C),.A2(FE_OFN289_g4679C),.A1(g554C));
AND2_X2 U_g5128C (.ZN(g5128C),.A2(FE_OFN352_g109C),.A1(I7048C));
AND2_X1 U_g4962C (.ZN(g4962C),.A2(g4467C),.A1(g1651C));
AND2_X1 U_g4358C (.ZN(g4358C),.A2(g3906C),.A1(g1209C));
AND2_X1 U_g8683C (.ZN(g8683C),.A2(g8549C),.A1(g4803C));
AND2_X1 U_g4506C (.ZN(g4506C),.A2(FE_OFN351_g3913C),.A1(g1113C));
AND2_X1 U_g6471C (.ZN(g6471C),.A2(g5878C),.A1(g5224C));
AND2_X1 U_g8778C (.ZN(g8778C),.A2(g1975C),.A1(g8688C));
AND2_X1 U_g11281C (.ZN(g11281C),.A2(g11203C),.A1(g4788C));
AND2_X1 U_g11146C (.ZN(g11146C),.A2(FE_OFN278_g10927C),.A1(g318C));
AND2_X1 U_g3904C (.ZN(g3904C),.A2(g627C),.A1(g2948C));
AND2_X1 U_g8075C (.ZN(g8075C),.A2(g7697C),.A1(g727C));
AND2_X1 U_g9829C (.ZN(g9829C),.A2(FE_OFN34_g9785C),.A1(g9723C));
AND3_X1 U_g8949C (.ZN(g8949C),.A3(g8828C),.A2(FE_OFN92_g2216C),.A1(g8255C));
AND2_X1 U_g7632C (.ZN(g7632C),.A2(g5420C),.A1(g7184C));
AND2_X1 U_g11290C (.ZN(g11290C),.A2(g4379C),.A1(g11246C));
AND2_X1 U_g6350C (.ZN(g6350C),.A2(FE_OFN346_g4381C),.A1(g5837C));
AND2_X1 U_g10599C (.ZN(g10599C),.A2(g4365C),.A1(g10448C));
AND2_X1 U_g5902C (.ZN(g5902C),.A2(g4977C),.A1(g2555C));
AND4_X1 U_I6337C (.ZN(I6337C),.A4(g2396C),.A3(g2407C),.A2(g2421C),.A1(g201C));
AND2_X2 U_g2276C (.ZN(g2276C),.A2(g1610C),.A1(g1765C));
AND2_X1 U_g6438C (.ZN(g6438C),.A2(g5013C),.A1(g5853C));
AND2_X1 U_g5512C (.ZN(g5512C),.A2(g4281C),.A1(g1660C));
AND2_X1 U_g5090C (.ZN(g5090C),.A2(FE_OFN299_g4457C),.A1(g1781C));
AND2_X1 U_g7719C (.ZN(g7719C),.A2(FE_OFN191_g6488C),.A1(g718C));
AND2_X1 U_g2561C (.ZN(g2561C),.A2(g741C),.A1(g742C));
AND2_X1 U_g3695C (.ZN(g3695C),.A2(FE_OFN292_g3015C),.A1(g1712C));
AND2_X1 U_g8603C (.ZN(g8603C),.A2(g8548C),.A1(g3983C));
AND2_X1 U_g8039C (.ZN(g8039C),.A2(FE_OFN305_g5151C),.A1(g7587C));
AND2_X1 U_g9610C (.ZN(g9610C),.A2(g9192C),.A1(g925C));
AND2_X1 U_g3536C (.ZN(g3536C),.A2(g3103C),.A1(g1289C));
AND2_X1 U_g5529C (.ZN(g5529C),.A2(FE_OFN310_g4336C),.A1(g2257C));
AND2_X1 U_g5148C (.ZN(g5148C),.A2(g4671C),.A1(g1107C));
AND2_X1 U_g9124C (.ZN(g9124C),.A2(FE_OFN325_g18C),.A1(g8881C));
AND2_X1 U_g9324C (.ZN(g9324C),.A2(FE_OFN275_g48C),.A1(g8879C));
AND2_X1 U_g4559C (.ZN(g4559C),.A2(FE_OFN137_g3829C),.A1(g2034C));
AND2_X1 U_g10561C (.ZN(g10561C),.A2(FE_OFN370_g4525C),.A1(g10549C));
AND2_X1 U_g5698C (.ZN(g5698C),.A2(FE_OFN315_g5117C),.A1(g1571C));
AND2_X1 U_g11226C (.ZN(g11226C),.A2(g11060C),.A1(g461C));
AND2_X1 U_g10295C (.ZN(g10295C),.A2(g9995C),.A1(FE_OFN79_g8700C));
AND2_X1 U_g5260C (.ZN(g5260C),.A2(FE_OFN288_g4263C),.A1(g1092C));
AND2_X1 U_g10680C (.ZN(g10680C),.A2(FE_OFN102_g3586C),.A1(g10564C));
AND2_X1 U_g6822C (.ZN(g6822C),.A2(FE_OFN178_g5354C),.A1(g231C));
AND2_X1 U_g4905C (.ZN(g4905C),.A2(g4243C),.A1(g1853C));
AND2_X1 U_g11551C (.ZN(g11551C),.A2(FE_OFN119_g3015C),.A1(g11538C));
AND2_X1 U_g3047C (.ZN(g3047C),.A2(g2306C),.A1(g1227C));
AND2_X1 U_g9849C (.ZN(g9849C),.A2(g9764C),.A1(g293C));
AND2_X1 U_g5279C (.ZN(g5279C),.A2(FE_OFN299_g4457C),.A1(g1766C));
AND2_X1 U_g8404C (.ZN(g8404C),.A2(g8146C),.A1(g686C));
AND2_X1 U_g5720C (.ZN(g5720C),.A2(FE_OFN168_g5361C),.A1(g170C));
AND2_X1 U_g5318C (.ZN(g5318C),.A2(g1857C),.A1(FE_OFN223_g4401C));
AND2_X1 U_g11376C (.ZN(g11376C),.A2(g4285C),.A1(g11318C));
AND2_X1 U_g11297C (.ZN(g11297C),.A2(g11243C),.A1(g4565C));
AND2_X1 U_g9898C (.ZN(g9898C),.A2(g9367C),.A1(g9710C));
OR2_X1 U_g6895C (.ZN(g6895C),.A2(g4875C),.A1(g6776C));
OR2_X1 U_g7189C (.ZN(g7189C),.A2(I9717C),.A1(g6632C));
OR2_X1 U_g9510C (.ZN(g9510C),.A2(g9111C),.A1(FE_OFN44_g9125C));
OR2_X1 U_g7297C (.ZN(g7297C),.A2(g6323C),.A1(g7132C));
OR2_X1 U_g9088C (.ZN(g9088C),.A2(g8233C),.A1(g8927C));
OR2_X1 U_g9923C (.ZN(g9923C),.A2(g9707C),.A1(g9865C));
OR2_X1 U_g6485C (.ZN(g6485C),.A2(g5067C),.A1(g5848C));
OR2_X1 U_g8771C (.ZN(g8771C),.A2(g8652C),.A1(g5483C));
OR2_X1 U_g5813C (.ZN(g5813C),.A2(g4869C),.A1(g5617C));
OR2_X1 U_g7963C (.ZN(g7963C),.A2(g7182C),.A1(FE_OFN334_g7045C));
OR2_X1 U_g10643C (.ZN(g10643C),.A2(g7736C),.A1(g10624C));
OR3_X1 U_g9886C (.ZN(g9886C),.A3(g9759C),.A2(g9592C),.A1(g9607C));
OR3_X1 U_g9951C (.ZN(g9951C),.A3(g9803C),.A2(g9899C),.A1(g9902C));
OR2_X1 U_g11625C (.ZN(g11625C),.A2(g11597C),.A1(g6535C));
OR2_X1 U_g8945C (.ZN(g8945C),.A2(FE_OFN332_g8748C),.A1(g8801C));
OR2_X1 U_g10489C (.ZN(g10489C),.A2(g10367C),.A1(g4456C));
OR2_X1 U_g10559C (.ZN(g10559C),.A2(g10512C),.A1(g4141C));
OR2_X1 U_g10558C (.ZN(g10558C),.A2(g10510C),.A1(g4126C));
OR2_X1 U_g11338C (.ZN(g11338C),.A2(g11178C),.A1(g11283C));
OR2_X1 U_g8435C (.ZN(g8435C),.A2(g8075C),.A1(g8403C));
OR2_X1 U_g10544C (.ZN(g10544C),.A2(g10495C),.A1(g4271C));
OR2_X1 U_g6911C (.ZN(g6911C),.A2(g5681C),.A1(g6342C));
OR2_X1 U_g10865C (.ZN(g10865C),.A2(g10752C),.A1(g5538C));
OR2_X1 U_g3698C (.ZN(g3698C),.A2(g869C),.A1(g3121C));
OR2_X1 U_g8214C (.ZN(g8214C),.A2(g7682C),.A1(g7472C));
OR2_X1 U_g6124C (.ZN(g6124C),.A2(g5188C),.A1(g5181C));
OR2_X1 U_g6469C (.ZN(g6469C),.A2(g4959C),.A1(g5698C));
OR2_X1 U_g5587C (.ZN(g5587C),.A2(g3904C),.A1(g4714C));
OR2_X1 U_g6177C (.ZN(g6177C),.A2(g4712C),.A1(g5444C));
OR2_X1 U_g9891C (.ZN(g9891C),.A2(g9760C),.A1(FE_OFN33_g9454C));
OR2_X1 U_g9913C (.ZN(g9913C),.A2(g9691C),.A1(g9849C));
OR4_X1 U_I5600C (.ZN(I5600C),.A4(g481C),.A3(g486C),.A2(g491C),.A1(g496C));
OR2_X1 U_g11257C (.ZN(g11257C),.A2(g11019C),.A1(g11234C));
OR2_X1 U_g8236C (.ZN(g8236C),.A2(g7680C),.A1(g7526C));
OR2_X1 U_g7385C (.ZN(g7385C),.A2(g6746C),.A1(g7235C));
OR2_X1 U_g6898C (.ZN(g6898C),.A2(g4881C),.A1(g6790C));
OR2_X1 U_g6900C (.ZN(g6900C),.A2(g6246C),.A1(g6787C));
OR2_X1 U_g4264C (.ZN(g4264C),.A2(g4053C),.A1(g4048C));
OR3_X1 U_g9726C (.ZN(g9726C),.A3(g9426C),.A2(g9420C),.A1(g9411C));
OR2_X1 U_g6088C (.ZN(g6088C),.A2(g4522C),.A1(g5260C));
OR2_X1 U_g6923C (.ZN(g6923C),.A2(g5695C),.A1(g6353C));
OR2_X1 U_g8194C (.ZN(g8194C),.A2(g7940C),.A1(g5168C));
OR3_X1 U_g9676C (.ZN(g9676C),.A3(FE_OFN62_g9274C),.A2(FE_OFN72_g9292C),.A1(g9454C));
OR2_X1 U_g11256C (.ZN(g11256C),.A2(g11018C),.A1(g11186C));
OR2_X1 U_g3860C (.ZN(g3860C),.A2(g2167C),.A1(g3107C));
OR2_X1 U_g11280C (.ZN(g11280C),.A2(g11153C),.A1(g11254C));
OR4_X1 U_g9727C (.ZN(g9727C),.A4(I14866C),.A3(g9391C),.A2(g9663C),.A1(g9650C));
OR2_X1 U_g4997C (.ZN(g4997C),.A2(g4584C),.A1(g4581C));
OR2_X1 U_g11624C (.ZN(g11624C),.A2(g11571C),.A1(g11595C));
OR2_X1 U_g11300C (.ZN(g11300C),.A2(g11091C),.A1(g11213C));
OR2_X1 U_g4238C (.ZN(g4238C),.A2(g4007C),.A1(g3999C));
OR2_X1 U_g8814C (.ZN(g8814C),.A2(g8728C),.A1(g7945C));
OR2_X1 U_g10401C (.ZN(g10401C),.A2(g10291C),.A1(g9317C));
OR2_X1 U_g8773C (.ZN(g8773C),.A2(g8653C),.A1(g5491C));
OR2_X1 U_g11231C (.ZN(g11231C),.A2(g11013C),.A1(g11156C));
OR2_X1 U_g10864C (.ZN(g10864C),.A2(g10751C),.A1(g5532C));
OR2_X1 U_g9624C (.ZN(g9624C),.A2(g9313C),.A1(g9316C));
OR3_X1 U_g9953C (.ZN(g9953C),.A3(g9803C),.A2(g9939C),.A1(g9945C));
OR2_X1 U_g6122C (.ZN(g6122C),.A2(g5180C),.A1(g5172C));
OR2_X1 U_g6465C (.ZN(g6465C),.A2(g5041C),.A1(g5825C));
OR2_X1 U_g6934C (.ZN(g6934C),.A2(g5720C),.A1(g6363C));
OR2_X1 U_g7664C (.ZN(g7664C),.A2(FE_OFN350_g3121C),.A1(g6855C));
OR2_X1 U_g7246C (.ZN(g7246C),.A2(g6003C),.A1(g6465C));
OR2_X1 U_g7203C (.ZN(g7203C),.A2(g6058C),.A1(g6640C));
OR2_X1 U_g6096C (.ZN(g6096C),.A2(g4542C),.A1(g5268C));
OR2_X1 U_g9747C (.ZN(g9747C),.A2(g9509C),.A1(g9173C));
OR2_X1 U_g11314C (.ZN(g11314C),.A2(g11102C),.A1(g11224C));
OR2_X1 U_g10733C (.ZN(g10733C),.A2(g10679C),.A1(g5227C));
OR2_X1 U_g8921C (.ZN(g8921C),.A2(g8748C),.A1(g8827C));
OR4_X1 U_I15054C (.ZN(I15054C),.A4(FE_OFN35_g9785C),.A3(FE_OFN61_g9624C),.A2(FE_OFN32_g9454C),.A1(FE_OFN90_I11360C));
OR2_X1 U_g11269C (.ZN(g11269C),.A2(g11031C),.A1(g11196C));
OR2_X1 U_g5555C (.ZN(g5555C),.A2(g4397C),.A1(g4389C));
OR2_X1 U_g11268C (.ZN(g11268C),.A2(g11030C),.A1(g11194C));
OR2_X1 U_g10485C (.ZN(g10485C),.A2(g10363C),.A1(g9317C));
OR2_X1 U_g10555C (.ZN(g10555C),.A2(g10504C),.A1(g4103C));
OR2_X1 U_g6481C (.ZN(g6481C),.A2(g4972C),.A1(g5722C));
OR2_X1 U_g10712C (.ZN(g10712C),.A2(g9097C),.A1(g10662C));
OR2_X1 U_g11335C (.ZN(g11335C),.A2(g11175C),.A1(g11279C));
OR2_X1 U_g8249C (.ZN(g8249C),.A2(g7710C),.A1(g8018C));
OR2_X1 U_g7638C (.ZN(g7638C),.A2(FE_OFN195_g6488C),.A1(g7265C));
OR2_X1 U_g10567C (.ZN(g10567C),.A2(g7378C),.A1(g10514C));
OR2_X1 U_g11487C (.ZN(g11487C),.A2(g11464C),.A1(g6662C));
OR4_X1 U_I15210C (.ZN(I15210C),.A4(g9882C),.A3(g9852C),.A2(g9964C),.A1(g9839C));
OR4_X1 U_I5805C (.ZN(I5805C),.A4(g2088C),.A3(g2096C),.A2(g2099C),.A1(g2102C));
OR2_X1 U_g8941C (.ZN(g8941C),.A2(FE_OFN332_g8748C),.A1(g8796C));
OR2_X1 U_g11443C (.ZN(g11443C),.A2(g11407C),.A1(g7130C));
OR2_X1 U_g4231C (.ZN(g4231C),.A2(g3998C),.A1(g3991C));
OR2_X1 U_g11278C (.ZN(g11278C),.A2(g11150C),.A1(g11253C));
OR2_X1 U_g11286C (.ZN(g11286C),.A2(g11209C),.A1(g10670C));
OR2_X1 U_g8431C (.ZN(g8431C),.A2(g8071C),.A1(g8387C));
OR2_X1 U_g7133C (.ZN(g7133C),.A2(I6273C),.A1(g6616C));
OR2_X1 U_g11306C (.ZN(g11306C),.A2(g11095C),.A1(g11216C));
OR2_X1 U_g8252C (.ZN(g8252C),.A2(g7679C),.A1(g7988C));
OR2_X1 U_g8812C (.ZN(g8812C),.A2(g8724C),.A1(g7939C));
OR2_X1 U_g7846C (.ZN(g7846C),.A2(g7241C),.A1(g7722C));
OR2_X1 U_g3875C (.ZN(g3875C),.A2(g12C),.A1(g3275C));
OR2_X1 U_g5996C (.ZN(g5996C),.A2(g3383C),.A1(g5473C));
OR2_X1 U_g6592C (.ZN(g6592C),.A2(g5882C),.A1(g5100C));
OR2_X1 U_g8286C (.ZN(g8286C),.A2(g7823C),.A1(g8107C));
OR2_X1 U_g10501C (.ZN(g10501C),.A2(g10445C),.A1(g4161C));
OR2_X1 U_g10728C (.ZN(g10728C),.A2(g10642C),.A1(g4973C));
OR2_X1 U_g8270C (.ZN(g8270C),.A2(g3434C),.A1(g7894C));
OR2_X1 U_g7290C (.ZN(g7290C),.A2(g6316C),.A1(g7046C));
OR2_X1 U_g6068C (.ZN(g6068C),.A2(g4497C),.A1(g5220C));
OR2_X1 U_g6468C (.ZN(g6468C),.A2(g4950C),.A1(g5690C));
OR2_X1 U_g11217C (.ZN(g11217C),.A2(g11005C),.A1(g11144C));
OR2_X1 U_g11478C (.ZN(g11478C),.A2(g11455C),.A1(g6532C));
OR4_X2 U_g9536C (.ZN(g9536C),.A4(g9324C),.A3(g9328C),.A2(g9331C),.A1(g9335C));
OR2_X1 U_g5981C (.ZN(g5981C),.A2(g4383C),.A1(g5074C));
OR2_X1 U_g11486C (.ZN(g11486C),.A2(g11463C),.A1(g6654C));
OR2_X1 U_g8377C (.ZN(g8377C),.A2(g7958C),.A1(g8185C));
OR2_X1 U_g8206C (.ZN(g8206C),.A2(g7683C),.A1(g7459C));
OR2_X1 U_g11580C (.ZN(g11580C),.A2(g11544C),.A1(g11413C));
OR2_X1 U_g8287C (.ZN(g8287C),.A2(g7824C),.A1(g8117C));
OR2_X1 U_g11223C (.ZN(g11223C),.A2(g11008C),.A1(g11147C));
OR2_X1 U_g9522C (.ZN(g9522C),.A2(FE_OFN44_g9125C),.A1(g9173C));
OR2_X1 U_g8199C (.ZN(g8199C),.A2(g7444C),.A1(g7902C));
OR2_X1 U_g5802C (.ZN(g5802C),.A2(g4837C),.A1(g5601C));
OR2_X1 U_g11321C (.ZN(g11321C),.A2(g11105C),.A1(g11230C));
OR2_X1 U_g6524C (.ZN(g6524C),.A2(g4996C),.A1(g5746C));
OR2_X1 U_g10664C (.ZN(g10664C),.A2(g10582C),.A1(g10240C));
OR2_X1 U_g7257C (.ZN(g7257C),.A2(g4725C),.A1(g6701C));
OR2_X1 U_g7301C (.ZN(g7301C),.A2(g6327C),.A1(g7140C));
OR2_X1 U_g10484C (.ZN(g10484C),.A2(g10400C),.A1(g9317C));
OR2_X1 U_g10554C (.ZN(g10554C),.A2(g10503C),.A1(g4097C));
OR2_X1 U_g8259C (.ZN(g8259C),.A2(g7719C),.A1(g8028C));
OR2_X1 U_g11334C (.ZN(g11334C),.A2(g11174C),.A1(g11277C));
OR2_X1 U_g8819C (.ZN(g8819C),.A2(g8734C),.A1(g7957C));
OR2_X1 U_g8923C (.ZN(g8923C),.A2(FE_OFN329_g8763C),.A1(g8846C));
OR2_X2 U_g8488C (.ZN(g8488C),.A2(g8390C),.A1(FE_OFN204_g3664C));
OR2_X1 U_g7441C (.ZN(g7441C),.A2(g5867C),.A1(g7271C));
OR2_X1 U_g6026C (.ZN(g6026C),.A2(g3970C),.A1(g5507C));
OR2_X1 U_g10799C (.ZN(g10799C),.A2(g10769C),.A1(g6225C));
OR2_X1 U_g10798C (.ZN(g10798C),.A2(g10768C),.A1(g6217C));
OR2_X1 U_g10805C (.ZN(g10805C),.A2(g10760C),.A1(g10759C));
OR2_X1 U_g10732C (.ZN(g10732C),.A2(g10661C),.A1(g4358C));
OR2_X1 U_g6061C (.ZN(g6061C),.A2(g4C),.A1(g5204C));
OR2_X1 U_g9512C (.ZN(g9512C),.A2(g9125C),.A1(g9151C));
OR2_X1 U_g10013C (.ZN(g10013C),.A2(I15215C),.A1(I15214C));
OR2_X1 U_g8806C (.ZN(g8806C),.A2(g8718C),.A1(g7931C));
OR2_X1 U_g8943C (.ZN(g8943C),.A2(FE_OFN332_g8748C),.A1(g8837C));
OR2_X1 U_g11293C (.ZN(g11293C),.A2(g10818C),.A1(g11211C));
OR2_X1 U_g11265C (.ZN(g11265C),.A2(g11027C),.A1(g11189C));
OR2_X1 U_g8887C (.ZN(g8887C),.A2(FE_OFN329_g8763C),.A1(g8842C));
OR2_X1 U_g5838C (.ZN(g5838C),.A2(g3974C),.A1(g5612C));
OR2_X1 U_g6514C (.ZN(g6514C),.A2(g4992C),.A1(g5738C));
OR2_X1 U_g8322C (.ZN(g8322C),.A2(g6891C),.A1(g8136C));
OR2_X1 U_g8230C (.ZN(g8230C),.A2(g7686C),.A1(g7515C));
OR2_X1 U_g5809C (.ZN(g5809C),.A2(g4865C),.A1(g5611C));
OR2_X1 U_g8433C (.ZN(g8433C),.A2(g8073C),.A1(g8399C));
OR2_X1 U_g11579C (.ZN(g11579C),.A2(g11551C),.A1(g5123C));
OR2_X1 U_g10771C (.ZN(g10771C),.A2(g10684C),.A1(g5533C));
OR2_X1 U_g11615C (.ZN(g11615C),.A2(g11592C),.A1(g11601C));
OR2_X1 U_g9367C (.ZN(g9367C),.A2(g9331C),.A1(g9335C));
OR3_X1 U_g9872C (.ZN(g9872C),.A3(g9759C),.A2(g9594C),.A1(g9617C));
OR2_X1 U_g6522C (.ZN(g6522C),.A2(g4994C),.A1(g5744C));
OR2_X1 U_g8266C (.ZN(g8266C),.A2(g3412C),.A1(g7885C));
OR2_X1 U_g10414C (.ZN(g10414C),.A2(g9291C),.A1(g10300C));
OR2_X1 U_g11275C (.ZN(g11275C),.A2(g11148C),.A1(g11248C));
OR2_X1 U_g11430C (.ZN(g11430C),.A2(g4006C),.A1(g11387C));
OR2_X1 U_g8248C (.ZN(g8248C),.A2(g7707C),.A1(g8014C));
OR2_X1 U_g8815C (.ZN(g8815C),.A2(g8730C),.A1(g7948C));
OR2_X1 U_g7183C (.ZN(g7183C),.A2(I9717C),.A1(g6623C));
OR2_X1 U_g5983C (.ZN(g5983C),.A2(g4392C),.A1(g5084C));
OR2_X1 U_g8154C (.ZN(g8154C),.A2(g6879C),.A1(g7891C));
OR2_X1 U_g6537C (.ZN(g6537C),.A2(g5005C),.A1(g5781C));
OR2_X1 U_g4309C (.ZN(g4309C),.A2(g4079C),.A1(g4069C));
OR2_X1 U_g10725C (.ZN(g10725C),.A2(g10634C),.A1(g4962C));
OR2_X1 U_g6243C (.ZN(g6243C),.A2(g4144C),.A1(g5537C));
OR4_X1 U_I6351C (.ZN(I6351C),.A4(g2372C),.A3(g2380C),.A2(g2389C),.A1(g2405C));
OR3_X1 U_g9519C (.ZN(g9519C),.A3(FE_OFN44_g9125C),.A2(g9151C),.A1(g9173C));
OR2_X1 U_g9740C (.ZN(g9740C),.A2(g9505C),.A1(g9418C));
OR2_X1 U_g8267C (.ZN(g8267C),.A2(g3422C),.A1(g7889C));
OR3_X1 U_g10744C (.ZN(g10744C),.A3(I16427C),.A2(g10668C),.A1(g10381C));
OR2_X1 U_g6542C (.ZN(g6542C),.A2(g5010C),.A1(g5789C));
OR2_X1 U_g7303C (.ZN(g7303C),.A2(g6329C),.A1(g7145C));
OR2_X1 U_g10652C (.ZN(g10652C),.A2(g7743C),.A1(g10627C));
OR2_X1 U_g5036C (.ZN(g5036C),.A2(g4162C),.A1(g4871C));
OR2_X1 U_g7240C (.ZN(g7240C),.A2(g6095C),.A1(g6687C));
OR2_X1 U_g8221C (.ZN(g8221C),.A2(g7688C),.A1(g7496C));
OR2_X1 U_g6902C (.ZN(g6902C),.A2(g4223C),.A1(g6794C));
OR2_X1 U_g10500C (.ZN(g10500C),.A2(g10442C),.A1(g4157C));
OR2_X1 U_g4052C (.ZN(g4052C),.A2(g2515C),.A1(g2862C));
OR4_X1 U_I14858C (.ZN(I14858C),.A4(g9602C),.A3(g9610C),.A2(g9595C),.A1(g9585C));
OR2_X1 U_g6529C (.ZN(g6529C),.A2(g5000C),.A1(g5757C));
OR2_X1 U_g11264C (.ZN(g11264C),.A2(g11026C),.A1(g11188C));
OR4_X1 U_I15209C (.ZN(I15209C),.A4(g9830C),.A3(g9934C),.A2(g9905C),.A1(g8169C));
OR2_X1 U_g8241C (.ZN(g8241C),.A2(g7684C),.A1(g7536C));
OR2_X1 U_g10795C (.ZN(g10795C),.A2(g10764C),.A1(g6199C));
OR2_X1 U_g11607C (.ZN(g11607C),.A2(g11557C),.A1(g11586C));
OR2_X1 U_g8644C (.ZN(g8644C),.A2(g8464C),.A1(g8123C));
OR3_X1 U_g4682C (.ZN(g4682C),.A3(g1570C),.A2(g3348C),.A1(g3563C));
OR2_X1 U_g8818C (.ZN(g8818C),.A2(g8733C),.A1(g7955C));
OR2_X1 U_g2984C (.ZN(g2984C),.A2(g2522C),.A1(g2528C));
OR2_X1 U_g9931C (.ZN(g9931C),.A2(g9900C),.A1(g8931C));
OR2_X1 U_g3414C (.ZN(g3414C),.A2(g2917C),.A1(g2911C));
OR2_X1 U_g9515C (.ZN(g9515C),.A2(g9151C),.A1(g9173C));
OR2_X1 U_g10724C (.ZN(g10724C),.A2(g10672C),.A1(g10312C));
OR2_X1 U_g7294C (.ZN(g7294C),.A2(g6320C),.A1(g7068C));
OR2_X1 U_g5189C (.ZN(g5189C),.A2(FE_OFN292_g3015C),.A1(g4345C));
OR2_X1 U_g8614C (.ZN(g8614C),.A2(g8510C),.A1(g8365C));
OR2_X1 U_g3513C (.ZN(g3513C),.A2(g2180C),.A1(g3118C));
OR2_X1 U_g6909C (.ZN(g6909C),.A2(g5309C),.A1(g6346C));
OR4_X1 U_I5571C (.ZN(I5571C),.A4(g426C),.A3(g386C),.A2(g391C),.A1(g396C));
OR2_X1 U_g4283C (.ZN(g4283C),.A2(g4063C),.A1(g4059C));
OR2_X1 U_g8939C (.ZN(g8939C),.A2(FE_OFN332_g8748C),.A1(g8791C));
OR2_X1 U_g2514C (.ZN(g2514C),.A2(I5600C),.A1(I5599C));
OR2_X1 U_g11327C (.ZN(g11327C),.A2(g11167C),.A1(g11297C));
OR2_X1 U_g8187C (.ZN(g8187C),.A2(g7677C),.A1(g7542C));
OR2_X1 U_g11606C (.ZN(g11606C),.A2(g11556C),.A1(g11585C));
OR2_X1 U_g11303C (.ZN(g11303C),.A2(g11092C),.A1(g11214C));
OR2_X1 U_g5309C (.ZN(g5309C),.A2(g4401C),.A1(FE_OFN204_g3664C));
OR2_X1 U_g8200C (.ZN(g8200C),.A2(g7685C),.A1(g7535C));
OR3_X1 U_g2522C (.ZN(g2522C),.A3(I5629C),.A2(g829C),.A1(g833C));
OR4_X1 U_g2315C (.ZN(g2315C),.A4(I5363C),.A3(g1113C),.A2(g1166C),.A1(g1163C));
OR2_X1 U_g6506C (.ZN(g6506C),.A2(g4989C),.A1(g5731C));
OR2_X1 U_g10649C (.ZN(g10649C),.A2(g7741C),.A1(g10626C));
OR2_X1 U_g8159C (.ZN(g8159C),.A2(g6886C),.A1(g7895C));
OR2_X1 U_g7626C (.ZN(g7626C),.A2(g3440C),.A1(g7060C));
OR2_X1 U_g10770C (.ZN(g10770C),.A2(g10682C),.A1(g5525C));
OR2_X1 U_g11483C (.ZN(g11483C),.A2(g11460C),.A1(g6633C));
OR2_X1 U_g8811C (.ZN(g8811C),.A2(g8722C),.A1(g7935C));
OR3_X1 U_g8642C (.ZN(g8642C),.A3(g8465C),.A2(g31C),.A1(g30C));
OR2_X1 U_g6545C (.ZN(g6545C),.A2(g5025C),.A1(g5795C));
OR2_X1 U_g10767C (.ZN(g10767C),.A2(g10681C),.A1(g5500C));
OR2_X1 U_g11326C (.ZN(g11326C),.A2(g11166C),.A1(g11296C));
OR2_X1 U_g10898C (.ZN(g10898C),.A2(g10777C),.A1(g4220C));
OR2_X1 U_g11252C (.ZN(g11252C),.A2(g10969C),.A1(g11099C));
OR2_X1 U_g10719C (.ZN(g10719C),.A2(g10666C),.A1(g10303C));
OR2_X1 U_g4609C (.ZN(g4609C),.A2(g119C),.A1(g3275C));
OR2_X1 U_g6507C (.ZN(g6507C),.A2(g4990C),.A1(g5732C));
OR2_X1 U_g10718C (.ZN(g10718C),.A2(g10706C),.A1(g6238C));
OR2_X1 U_g10521C (.ZN(g10521C),.A2(I16149C),.A1(I16148C));
OR2_X1 U_g7075C (.ZN(g7075C),.A2(g6530C),.A1(g5104C));
OR2_X1 U_g7292C (.ZN(g7292C),.A2(g6318C),.A1(g7055C));
OR2_X1 U_g10861C (.ZN(g10861C),.A2(g10745C),.A1(g5523C));
OR2_X1 U_g8417C (.ZN(g8417C),.A2(g7721C),.A1(g8246C));
OR2_X1 U_g6515C (.ZN(g6515C),.A2(g4993C),.A1(g5739C));
OR4_X1 U_I14855C (.ZN(I14855C),.A4(g9596C),.A3(g9601C),.A2(g9593C),.A1(g9583C));
OR4_X1 U_I15205C (.ZN(I15205C),.A4(g9878C),.A3(g9850C),.A2(g9963C),.A1(g9838C));
OR4_X1 U_I15051C (.ZN(I15051C),.A4(FE_OFN35_g9785C),.A3(FE_OFN60_g9624C),.A2(g9673C),.A1(FE_OFN90_I11360C));
OR3_X1 U_g9724C (.ZN(g9724C),.A3(g9426C),.A2(g9419C),.A1(g9409C));
OR2_X1 U_g6528C (.ZN(g6528C),.A2(g4999C),.A1(g5756C));
OR2_X1 U_g8823C (.ZN(g8823C),.A2(g8693C),.A1(g8778C));
OR2_X1 U_g7503C (.ZN(g7503C),.A2(g6430C),.A1(g6887C));
OR2_X1 U_g8148C (.ZN(g8148C),.A2(g6872C),.A1(g7884C));
OR2_X1 U_g8649C (.ZN(g8649C),.A2(g3440C),.A1(g8499C));
OR2_X1 U_g3584C (.ZN(g3584C),.A2(g2516C),.A1(g2863C));
OR2_X1 U_g10776C (.ZN(g10776C),.A2(g10758C),.A1(g5544C));
OR3_X1 U_g9680C (.ZN(g9680C),.A3(FE_OFN62_g9274C),.A2(FE_OFN72_g9292C),.A1(FE_OFN32_g9454C));
OR2_X1 U_g10859C (.ZN(g10859C),.A2(g10742C),.A1(g5512C));
OR3_X1 U_I14866C (.ZN(I14866C),.A3(g9619C),.A2(g9609C),.A1(g9590C));
OR2_X1 U_g7299C (.ZN(g7299C),.A2(g6325C),.A1(g7138C));
OR2_X1 U_g10858C (.ZN(g10858C),.A2(g10741C),.A1(g5501C));
OR2_X1 U_g8193C (.ZN(g8193C),.A2(g7937C),.A1(g5145C));
OR3_X1 U_g9511C (.ZN(g9511C),.A3(g9111C),.A2(g9125C),.A1(g9151C));
OR2_X1 U_g7738C (.ZN(g7738C),.A2(g6738C),.A1(g7200C));
OR2_X1 U_g7244C (.ZN(g7244C),.A2(g4720C),.A1(g6699C));
OR2_X1 U_g3425C (.ZN(g3425C),.A2(g2910C),.A1(g2895C));
OR2_X1 U_g7478C (.ZN(g7478C),.A2(g6423C),.A1(g6884C));
OR3_X1 U_g9714C (.ZN(g9714C),.A3(g9654C),.A2(g9366C),.A1(g9664C));
OR2_X1 U_g10025C (.ZN(g10025C),.A2(I15225C),.A1(I15224C));
OR2_X1 U_g6908C (.ZN(g6908C),.A2(g4229C),.A1(g6345C));
OR2_X1 U_g5028C (.ZN(g5028C),.A2(g4128C),.A1(g4836C));
OR2_X1 U_g8253C (.ZN(g8253C),.A2(g7718C),.A1(g8023C));
OR2_X1 U_g8938C (.ZN(g8938C),.A2(FE_OFN332_g8748C),.A1(g8789C));
OR2_X1 U_g8813C (.ZN(g8813C),.A2(g8726C),.A1(g7943C));
OR2_X1 U_g9736C (.ZN(g9736C),.A2(g9423C),.A1(g9430C));
OR2_X1 U_g9968C (.ZN(g9968C),.A2(I15172C),.A1(I15171C));
OR2_X1 U_g8552C (.ZN(g8552C),.A2(g8388C),.A1(g8217C));
OR2_X1 U_g5910C (.ZN(g5910C),.A2(g4341C),.A1(g5023C));
OR2_X1 U_g11249C (.ZN(g11249C),.A2(g11143C),.A1(g6162C));
OR2_X1 U_g11482C (.ZN(g11482C),.A2(g11459C),.A1(g6628C));
OR4_X1 U_g9722C (.ZN(g9722C),.A4(I14855C),.A3(g9391C),.A2(g9643C),.A1(g9612C));
OR4_X1 U_I15204C (.ZN(I15204C),.A4(g9829C),.A3(g9933C),.A2(g9904C),.A1(g8168C));
OR2_X1 U_g7236C (.ZN(g7236C),.A2(g6092C),.A1(g6684C));
OR2_X1 U_g8645C (.ZN(g8645C),.A2(g8469C),.A1(g8127C));
OR2_X1 U_g11647C (.ZN(g11647C),.A2(g11637C),.A1(g6622C));
OR2_X1 U_g6777C (.ZN(g6777C),.A2(g48C),.A1(I9221C));
OR3_X1 U_g9737C (.ZN(g9737C),.A3(g9387C),.A2(g9658C),.A1(g9657C));
OR4_X1 U_I16149C (.ZN(I16149C),.A4(g10467C),.A3(g10468C),.A2(g10470C),.A1(g10472C));
OR2_X1 U_g11233C (.ZN(g11233C),.A2(g10946C),.A1(g11085C));
OR2_X1 U_g8607C (.ZN(g8607C),.A2(g8554C),.A1(g8406C));
OR4_X1 U_I16148C (.ZN(I16148C),.A4(g10474C),.A3(g10476C),.A2(g10384C),.A1(g10386C));
OR2_X1 U_g8158C (.ZN(g8158C),.A2(g6883C),.A1(g7893C));
OR2_X1 U_g5846C (.ZN(g5846C),.A2(g4236C),.A1(g4932C));
OR2_X1 U_g5396C (.ZN(g5396C),.A2(g3684C),.A1(g4481C));
OR2_X1 U_g5803C (.ZN(g5803C),.A2(g3383C),.A1(g5575C));
OR2_X1 U_g11331C (.ZN(g11331C),.A2(g11171C),.A1(g11272C));
OR2_X1 U_g7295C (.ZN(g7295C),.A2(g6321C),.A1(g7071C));
OR2_X1 U_g6541C (.ZN(g6541C),.A2(g5009C),.A1(g5788C));
OR2_X1 U_g8615C (.ZN(g8615C),.A2(g8557C),.A1(g8413C));
OR2_X1 U_g9926C (.ZN(g9926C),.A2(g9715C),.A1(g9868C));
OR2_X1 U_g9754C (.ZN(g9754C),.A2(g9511C),.A1(g9173C));
OR2_X1 U_g8284C (.ZN(g8284C),.A2(g7821C),.A1(g8102C));
OR2_X1 U_g2204C (.ZN(g2204C),.A2(g1394C),.A1(g1393C));
OR2_X1 U_g7471C (.ZN(g7471C),.A2(g6416C),.A1(g6880C));
OR2_X1 U_g7242C (.ZN(g7242C),.A2(g6098C),.A1(g6693C));
OR2_X1 U_g5847C (.ZN(g5847C),.A2(g3987C),.A1(g5626C));
OR2_X1 U_g6901C (.ZN(g6901C),.A2(g6247C),.A1(g6788C));
OR2_X1 U_g8559C (.ZN(g8559C),.A2(g3664C),.A1(g8380C));
OR3_X1 U_g9729C (.ZN(g9729C),.A3(g9387C),.A2(g9357C),.A1(g9618C));
OR2_X1 U_g10860C (.ZN(g10860C),.A2(g10743C),.A1(g5513C));
OR2_X1 U_g9927C (.ZN(g9927C),.A2(g9716C),.A1(g9869C));
OR2_X1 U_g10497C (.ZN(g10497C),.A2(g10396C),.A1(FE_OFN277_g48C));
OR4_X1 U_g9885C (.ZN(g9885C),.A4(g9759C),.A3(g9662C),.A2(g9598C),.A1(g9454C));
OR4_X1 U_g2528C (.ZN(g2528C),.A4(g849C),.A3(g853C),.A2(g857C),.A1(g861C));
OR2_X1 U_g11229C (.ZN(g11229C),.A2(g11012C),.A1(g11154C));
OR2_X1 U_g8973C (.ZN(g8973C),.A2(FE_OFN329_g8763C),.A1(g8821C));
OR2_X1 U_g10658C (.ZN(g10658C),.A2(g7674C),.A1(g10595C));
OR2_X1 U_g10339C (.ZN(g10339C),.A2(g9291C),.A1(g10232C));
OR4_X1 U_I5363C (.ZN(I5363C),.A4(g1160C),.A3(g1157C),.A2(g1153C),.A1(g1149C));
OR2_X1 U_g11310C (.ZN(g11310C),.A2(g11100C),.A1(g11220C));
OR2_X1 U_g6500C (.ZN(g6500C),.A2(g4986C),.A1(g5725C));
OR2_X1 U_g10855C (.ZN(g10855C),.A2(g10736C),.A1(g6075C));
OR2_X1 U_g9916C (.ZN(g9916C),.A2(g9694C),.A1(g9855C));
OR2_X1 U_g10411C (.ZN(g10411C),.A2(g9291C),.A1(g10299C));
OR2_X1 U_g11603C (.ZN(g11603C),.A2(g11553C),.A1(g11582C));
OR4_X1 U_I5357C (.ZN(I5357C),.A4(g1250C),.A3(g1255C),.A2(g1260C),.A1(g1265C));
OR2_X1 U_g6672C (.ZN(g6672C),.A2(g5259C),.A1(g5509C));
OR3_X1 U_g9873C (.ZN(g9873C),.A3(g9758C),.A2(g9599C),.A1(g9623C));
OR2_X1 U_g6523C (.ZN(g6523C),.A2(g4995C),.A1(g5745C));
OR2_X1 U_g10707C (.ZN(g10707C),.A2(g10686C),.A1(g5545C));
OR4_X1 U_I5626C (.ZN(I5626C),.A4(g534C),.A3(g530C),.A2(g525C),.A1(g521C));
OR2_X1 U_g9579C (.ZN(g9579C),.A2(g9030C),.A1(FE_OFN54_g9052C));
OR2_X1 U_g7298C (.ZN(g7298C),.A2(g6324C),.A1(g7136C));
OR2_X1 U_g6551C (.ZN(g6551C),.A2(g5031C),.A1(g5804C));
OR2_X1 U_g6099C (.ZN(g6099C),.A2(g4550C),.A1(g5273C));
OR2_X1 U_g8282C (.ZN(g8282C),.A2(g7819C),.A1(g8101C));
OR2_X1 U_g9917C (.ZN(g9917C),.A2(g9695C),.A1(g9856C));
OR4_X1 U_I15057C (.ZN(I15057C),.A4(FE_OFN35_g9785C),.A3(FE_OFN60_g9624C),.A2(g9680C),.A1(FE_OFN90_I11360C));
OR2_X1 U_g7219C (.ZN(g7219C),.A2(I9717C),.A1(g6661C));
OR2_X1 U_g10019C (.ZN(g10019C),.A2(I15220C),.A1(I15219C));
OR2_X1 U_g5857C (.ZN(g5857C),.A2(g4670C),.A1(g5418C));
OR4_X1 U_g9725C (.ZN(g9725C),.A4(I14862C),.A3(g9391C),.A2(g9659C),.A1(g9642C));
OR2_X1 U_g11298C (.ZN(g11298C),.A2(g11087C),.A1(g11212C));
OR2_X1 U_g10402C (.ZN(g10402C),.A2(g9291C),.A1(g10295C));
OR4_X1 U_g2521C (.ZN(g2521C),.A4(I5626C),.A3(g476C),.A2(g542C),.A1(g538C));
OR2_X1 U_g10866C (.ZN(g10866C),.A2(g10753C),.A1(g5539C));
OR2_X1 U_g6534C (.ZN(g6534C),.A2(g5003C),.A1(g5772C));
OR2_X1 U_g11232C (.ZN(g11232C),.A2(g11015C),.A1(g11158C));
OR3_X1 U_g9706C (.ZN(g9706C),.A3(g9591C),.A2(g9386C),.A1(g9644C));
OR2_X1 U_g10001C (.ZN(g10001C),.A2(I15205C),.A1(I15204C));
OR2_X1 U_g8776C (.ZN(g8776C),.A2(g8655C),.A1(g5510C));
OR2_X1 U_g7225C (.ZN(g7225C),.A2(g6079C),.A1(g6666C));
OR3_X1 U_g9888C (.ZN(g9888C),.A3(g9757C),.A2(g9608C),.A1(g9648C));
OR2_X1 U_g11261C (.ZN(g11261C),.A2(g11023C),.A1(g11238C));
OR3_X1 U_g9956C (.ZN(g9956C),.A3(g9815C),.A2(g9942C),.A1(g9948C));
OR2_X1 U_g10923C (.ZN(g10923C),.A2(g10715C),.A1(g10778C));
OR2_X1 U_g8264C (.ZN(g8264C),.A2(g3912C),.A1(g7879C));
OR2_X1 U_g6513C (.ZN(g6513C),.A2(g4991C),.A1(g5737C));
OR3_X1 U_I14835C (.ZN(I14835C),.A3(g9588C),.A2(g9645C),.A1(g9621C));
OR2_X1 U_g8641C (.ZN(g8641C),.A2(g8463C),.A1(g8120C));
OR3_X1 U_g5361C (.ZN(g5361C),.A3(g126C),.A2(g3348C),.A1(g4316C));
OR2_X1 U_g11316C (.ZN(g11316C),.A2(g11103C),.A1(g11226C));
OR4_X1 U_I16161C (.ZN(I16161C),.A4(g10475C),.A3(g10477C),.A2(g10478C),.A1(g10479C));
OR2_X1 U_g6916C (.ZN(g6916C),.A2(g5687C),.A1(g6348C));
OR2_X1 U_g8777C (.ZN(g8777C),.A2(g8659C),.A1(g5522C));
OR4_X1 U_g2353C (.ZN(g2353C),.A4(g1415C),.A3(g1411C),.A2(g1407C),.A1(g1403C));
OR2_X1 U_g7510C (.ZN(g7510C),.A2(g6730C),.A1(g7186C));
OR3_X1 U_g9957C (.ZN(g9957C),.A3(g9803C),.A2(g9943C),.A1(g9949C));
OR2_X1 U_g2744C (.ZN(g2744C),.A2(I5805C),.A1(I5804C));
OR2_X1 U_g7245C (.ZN(g7245C),.A2(g6102C),.A1(g6696C));
OR2_X1 U_g7291C (.ZN(g7291C),.A2(g6317C),.A1(g7050C));
OR2_X1 U_g8611C (.ZN(g8611C),.A2(g8556C),.A1(g8410C));
OR4_X1 U_I15199C (.ZN(I15199C),.A4(g9828C),.A3(g9932C),.A2(g9903C),.A1(g8167C));
OR2_X1 U_g10550C (.ZN(g10550C),.A2(g10450C),.A1(g4437C));
OR2_X1 U_g11330C (.ZN(g11330C),.A2(g11170C),.A1(g11304C));
OR2_X1 U_g10721C (.ZN(g10721C),.A2(g10669C),.A1(g10306C));
OR2_X1 U_g8153C (.ZN(g8153C),.A2(g6875C),.A1(g7888C));
OR2_X1 U_g10773C (.ZN(g10773C),.A2(g10685C),.A1(g5540C));
OR2_X1 U_g3688C (.ZN(g3688C),.A2(g868C),.A1(g3744C));
OR4_X1 U_I15225C (.ZN(I15225C),.A4(g9881C),.A3(g9859C),.A2(g9967C),.A1(g9842C));
OR2_X1 U_g6042C (.ZN(g6042C),.A2(g3987C),.A1(g5535C));
OR2_X1 U_g10655C (.ZN(g10655C),.A2(g7389C),.A1(g10561C));
OR2_X1 U_g11259C (.ZN(g11259C),.A2(g11021C),.A1(g11236C));
OR2_X1 U_g11225C (.ZN(g11225C),.A2(g11009C),.A1(g11149C));
OR2_X1 U_g5914C (.ZN(g5914C),.A2(g4343C),.A1(g5029C));
OR2_X1 U_g11258C (.ZN(g11258C),.A2(g11020C),.A1(g11235C));
OR2_X1 U_g6054C (.ZN(g6054C),.A2(g4483C),.A1(g5199C));
OR3_X1 U_g9728C (.ZN(g9728C),.A3(g9426C),.A2(g9422C),.A1(g9412C));
OR3_X1 U_g9730C (.ZN(g9730C),.A3(g9423C),.A2(g9425C),.A1(g9414C));
OR2_X1 U_g5820C (.ZN(g5820C),.A2(g3942C),.A1(g5595C));
OR3_X1 U_g8574C (.ZN(g8574C),.A3(g8465C),.A2(I11360C),.A1(g30C));
OR2_X1 U_g11602C (.ZN(g11602C),.A2(g11552C),.A1(g11581C));
OR2_X1 U_g10502C (.ZN(g10502C),.A2(g10503C),.A1(g4169C));
OR2_X1 U_g10557C (.ZN(g10557C),.A2(g10508C),.A1(g4123C));
OR4_X1 U_I15171C (.ZN(I15171C),.A4(g9835C),.A3(g9896C),.A2(g9909C),.A1(g8175C));
OR2_X1 U_g11337C (.ZN(g11337C),.A2(g11177C),.A1(g11282C));
OR2_X1 U_g7465C (.ZN(g7465C),.A2(g6410C),.A1(g6876C));
OR2_X1 U_g8262C (.ZN(g8262C),.A2(g7625C),.A1(g7970C));
OR2_X1 U_g8889C (.ZN(g8889C),.A2(FE_OFN329_g8763C),.A1(g8844C));
OR2_X1 U_g7096C (.ZN(g7096C),.A2(g5911C),.A1(g6544C));
OR2_X1 U_g5995C (.ZN(g5995C),.A2(g5099C),.A1(g5097C));
OR2_X1 U_g8285C (.ZN(g8285C),.A2(g7822C),.A1(g8104C));
OR2_X1 U_g10791C (.ZN(g10791C),.A2(g10762C),.A1(g6186C));
OR2_X1 U_g2499C (.ZN(g2499C),.A2(I5571C),.A1(I5570C));
OR2_X1 U_g6049C (.ZN(g6049C),.A2(g4670C),.A1(g5254C));
OR2_X1 U_g9920C (.ZN(g9920C),.A2(g9701C),.A1(g9860C));
OR2_X1 U_g10556C (.ZN(g10556C),.A2(g10506C),.A1(g4115C));
OR2_X1 U_g8643C (.ZN(g8643C),.A2(g8508C),.A1(g8364C));
OR2_X1 U_g5810C (.ZN(g5810C),.A2(g3912C),.A1(g5588C));
OR2_X1 U_g11336C (.ZN(g11336C),.A2(g11176C),.A1(g11281C));
OR2_X1 U_g8742C (.ZN(g8742C),.A2(g8598C),.A1(g8135C));
OR2_X1 U_g8926C (.ZN(g8926C),.A2(g8763C),.A1(g8848C));
OR2_X1 U_g7218C (.ZN(g7218C),.A2(g6070C),.A1(g6655C));
OR4_X1 U_I15224C (.ZN(I15224C),.A4(g9834C),.A3(g9937C),.A2(g9908C),.A1(g8174C));
OR2_X1 U_g7293C (.ZN(g7293C),.A2(g6319C),.A1(g7063C));
OR2_X1 U_g11288C (.ZN(g11288C),.A2(g11070C),.A1(g11204C));
OR2_X1 U_g10800C (.ZN(g10800C),.A2(g10772C),.A1(g6245C));
OR2_X1 U_g11308C (.ZN(g11308C),.A2(g11098C),.A1(g11218C));
OR2_X1 U_g8269C (.ZN(g8269C),.A2(g3429C),.A1(g7892C));
OR2_X1 U_g10417C (.ZN(g10417C),.A2(g9097C),.A1(g10301C));
OR2_X1 U_g10936C (.ZN(g10936C),.A2(g10808C),.A1(g5170C));
OR2_X1 U_g9388C (.ZN(g9388C),.A2(g9223C),.A1(g9240C));
OR2_X1 U_g6185C (.ZN(g6185C),.A2(g4715C),.A1(g5470C));
OR2_X1 U_g6470C (.ZN(g6470C),.A2(g4960C),.A1(g5699C));
OR2_X1 U_g6897C (.ZN(g6897C),.A2(g6240C),.A1(g6771C));
OR2_X1 U_g8885C (.ZN(g8885C),.A2(FE_OFN329_g8763C),.A1(g8841C));
OR2_X1 U_g11260C (.ZN(g11260C),.A2(g11022C),.A1(g11237C));
OR2_X1 U_g11488C (.ZN(g11488C),.A2(g11465C),.A1(g6671C));
OR2_X1 U_g6105C (.ZN(g6105C),.A2(g4559C),.A1(g5279C));
OR2_X1 U_g10807C (.ZN(g10807C),.A2(g10761C),.A1(g10701C));
OR2_X1 U_g10639C (.ZN(g10639C),.A2(g7734C),.A1(g10623C));
OR2_X1 U_g4556C (.ZN(g4556C),.A2(g1212C),.A1(g3536C));
OR2_X1 U_g8288C (.ZN(g8288C),.A2(g7825C),.A1(g8119C));
OR2_X1 U_g6755C (.ZN(g6755C),.A2(g5479C),.A1(g4934C));
OR3_X1 U_I14862C (.ZN(I14862C),.A3(g9611C),.A2(g9600C),.A1(g9587C));
OR4_X1 U_I16160C (.ZN(I16160C),.A4(g10481C),.A3(g10482C),.A2(g10392C),.A1(g10394C));
OR2_X1 U_g11610C (.ZN(g11610C),.A2(g11560C),.A1(g11589C));
OR4_X1 U_g9711C (.ZN(g9711C),.A4(g9589C),.A3(g9359C),.A2(g9390C),.A1(g9660C));
OR2_X1 U_g6045C (.ZN(g6045C),.A2(g3989C),.A1(g5541C));
OR2_X1 U_g11270C (.ZN(g11270C),.A2(g11032C),.A1(g11198C));
OR2_X1 U_g7258C (.ZN(g7258C),.A2(g5913C),.A1(g6549C));
OR2_X1 U_g6059C (.ZN(g6059C),.A2(g4489C),.A1(g5211C));
OR2_X1 U_g10007C (.ZN(g10007C),.A2(I15210C),.A1(I15209C));
OR2_X1 U_g11267C (.ZN(g11267C),.A2(g11029C),.A1(g11192C));
OR2_X1 U_g11294C (.ZN(g11294C),.A2(g11210C),.A1(g6576C));
OR3_X1 U_g9509C (.ZN(g9509C),.A3(g9111C),.A2(FE_OFN44_g9125C),.A1(g9151C));
OR2_X1 U_g7211C (.ZN(g7211C),.A2(g6067C),.A1(g6647C));
OR2_X1 U_g5404C (.ZN(g5404C),.A2(g3696C),.A1(g4487C));
OR2_X1 U_g4089C (.ZN(g4089C),.A2(I5254C),.A1(g1959C));
OR4_X1 U_I15219C (.ZN(I15219C),.A4(g9833C),.A3(g9936C),.A2(g9907C),.A1(g8172C));
OR2_X1 U_g11219C (.ZN(g11219C),.A2(g11006C),.A1(g11145C));
OR2_X1 U_g6015C (.ZN(g6015C),.A2(g3942C),.A1(g5497C));
OR2_X1 U_g10720C (.ZN(g10720C),.A2(g10667C),.A1(g10304C));
OR2_X1 U_g8265C (.ZN(g8265C),.A2(g4827C),.A1(g7881C));
OR2_X1 U_g5224C (.ZN(g5224C),.A2(g3512C),.A1(g4360C));
OR3_X1 U_g9700C (.ZN(g9700C),.A3(I14827C),.A2(g9667C),.A1(g9358C));
OR2_X1 U_g7106C (.ZN(g7106C),.A2(g5917C),.A1(g6554C));
OR2_X1 U_g8770C (.ZN(g8770C),.A2(g8651C),.A1(g5476C));
OR2_X1 U_g11201C (.ZN(g11201C),.A2(g11011C),.A1(g11152C));
OR3_X1 U_g9950C (.ZN(g9950C),.A3(g9803C),.A2(g9898C),.A1(g9901C));
OR4_X1 U_g9723C (.ZN(g9723C),.A4(I14858C),.A3(g9391C),.A2(g9652C),.A1(g9620C));
OR2_X1 U_g2309C (.ZN(g2309C),.A2(I5358C),.A1(I5357C));
OR2_X1 U_g11266C (.ZN(g11266C),.A2(g11028C),.A1(g11190C));
OR2_X1 U_g10727C (.ZN(g10727C),.A2(g10638C),.A1(g4969C));
OR2_X1 U_g10863C (.ZN(g10863C),.A2(g10750C),.A1(g5531C));
OR2_X1 U_g8429C (.ZN(g8429C),.A2(g8069C),.A1(g8385C));
OR2_X1 U_g9751C (.ZN(g9751C),.A2(g9510C),.A1(g9515C));
OR2_X1 U_g8281C (.ZN(g8281C),.A2(g7818C),.A1(g8097C));
OR2_X1 U_g6910C (.ZN(g6910C),.A2(g5680C),.A1(g6341C));
OR2_X1 U_g8639C (.ZN(g8639C),.A2(g8462C),.A1(g8118C));
OR3_X1 U_g9673C (.ZN(g9673C),.A3(g9274C),.A2(FE_OFN72_g9292C),.A1(g9454C));
OR2_X1 U_g11285C (.ZN(g11285C),.A2(g11161C),.A1(g11255C));
OR2_X1 U_g11305C (.ZN(g11305C),.A2(g11093C),.A1(g11215C));
OR4_X1 U_I15177C (.ZN(I15177C),.A4(g9876C),.A3(g9863C),.A2(g9960C),.A1(g9844C));
OR3_X1 U_g9734C (.ZN(g9734C),.A3(g9426C),.A2(g9428C),.A1(g9415C));
OR3_X1 U_I14827C (.ZN(I14827C),.A3(g9584C),.A2(g9614C),.A1(g9603C));
OR2_X1 U_g5824C (.ZN(g5824C),.A2(g4839C),.A1(g5602C));
OR2_X1 U_g8715C (.ZN(g8715C),.A2(g8687C),.A1(g8416C));
OR2_X1 U_g5762C (.ZN(g5762C),.A2(g5186C),.A1(g5178C));
OR2_X1 U_g6538C (.ZN(g6538C),.A2(g5006C),.A1(g5782C));
OR2_X1 U_g5590C (.ZN(g5590C),.A2(g4723C),.A1(g4718C));
OR2_X1 U_g10726C (.ZN(g10726C),.A2(g10673C),.A1(g10316C));
OR2_X1 U_g3120C (.ZN(g3120C),.A2(I6351C),.A1(I6350C));
OR3_X2 U_g4640C (.ZN(g4640C),.A3(g1527C),.A2(g3563C),.A1(g3348C));
OR2_X1 U_g6093C (.ZN(g6093C),.A2(g4534C),.A1(g5264C));
OR2_X1 U_g8162C (.ZN(g8162C),.A2(g6889C),.A1(g7898C));
OR2_X1 U_g8268C (.ZN(g8268C),.A2(g7613C),.A1(g7962C));
OR2_X1 U_g9569C (.ZN(g9569C),.A2(FE_OFN49_g9030C),.A1(FE_OFN54_g9052C));
OR2_X1 U_g11485C (.ZN(g11485C),.A2(g11462C),.A1(g6646C));
OR2_X1 U_g10797C (.ZN(g10797C),.A2(g10766C),.A1(g6206C));
OR3_X1 U_I14779C (.ZN(I14779C),.A3(g9192C),.A2(g9205C),.A1(g8995C));
OR2_X1 U_g10408C (.ZN(g10408C),.A2(g9097C),.A1(g10298C));
OR2_X1 U_g10635C (.ZN(g10635C),.A2(g7732C),.A1(g10622C));
OR2_X1 U_g2305C (.ZN(g2305C),.A2(I5352C),.A1(I5351C));
OR4_X1 U_I15176C (.ZN(I15176C),.A4(g9836C),.A3(g9897C),.A2(g9908C),.A1(g8176C));
OR2_X1 U_g3435C (.ZN(g3435C),.A2(g2950C),.A1(g2945C));
OR2_X1 U_g9924C (.ZN(g9924C),.A2(g9709C),.A1(g9866C));
OR2_X1 U_g10711C (.ZN(g10711C),.A2(g10690C),.A1(g5547C));
OR2_X1 U_g5814C (.ZN(g5814C),.A2(g4827C),.A1(g5591C));
OR2_X1 U_g5038C (.ZN(g5038C),.A2(g4884C),.A1(g4878C));
OR4_X1 U_I15215C (.ZN(I15215C),.A4(g9879C),.A3(g9854C),.A2(g9965C),.A1(g9840C));
OR2_X1 U_g8226C (.ZN(g8226C),.A2(g7681C),.A1(g7504C));
OR2_X1 U_g7367C (.ZN(g7367C),.A2(g6744C),.A1(g7224C));
OR2_X1 U_g7457C (.ZN(g7457C),.A2(g6404C),.A1(g6873C));
OR2_X1 U_g5229C (.ZN(g5229C),.A2(g3516C),.A1(g4364C));
OR2_X1 U_g5993C (.ZN(g5993C),.A2(g4400C),.A1(g5090C));
OR2_X1 U_g8283C (.ZN(g8283C),.A2(g7820C),.A1(g8098C));
OR2_X1 U_g7971C (.ZN(g7971C),.A2(g7549C),.A1(g5110C));
OR2_X1 U_g8602C (.ZN(g8602C),.A2(g8550C),.A1(g8401C));
OR2_X1 U_g8920C (.ZN(g8920C),.A2(FE_OFN329_g8763C),.A1(g8845C));
OR2_X1 U_g10663C (.ZN(g10663C),.A2(g10581C),.A1(g10237C));
OR2_X1 U_g6074C (.ZN(g6074C),.A2(g1C),.A1(g5349C));
OR2_X1 U_g8261C (.ZN(g8261C),.A2(g3383C),.A1(g7876C));
OR2_X1 U_g10862C (.ZN(g10862C),.A2(g10746C),.A1(g5524C));
OR2_X1 U_g5837C (.ZN(g5837C),.A2(g4224C),.A1(g5640C));
OR2_X1 U_g11333C (.ZN(g11333C),.A2(g11173C),.A1(g11274C));
OR2_X1 U_g6080C (.ZN(g6080C),.A2(g4512C),.A1(g5249C));
OR2_X1 U_g6480C (.ZN(g6480C),.A2(g4971C),.A1(g5721C));
OR2_X1 U_g7740C (.ZN(g7740C),.A2(g6741C),.A1(g7209C));
OR2_X2 U_g10702C (.ZN(g10702C),.A2(g2984C),.A1(g10562C));
OR3_X1 U_g9697C (.ZN(g9697C),.A3(I14822C),.A2(g9606C),.A1(g9665C));
OR2_X1 U_g8203C (.ZN(g8203C),.A2(g7696C),.A1(g7453C));
OR2_X1 U_g9914C (.ZN(g9914C),.A2(g9692C),.A1(g9851C));
OR2_X1 U_g10564C (.ZN(g10564C),.A2(g7368C),.A1(g10560C));
OR2_X1 U_g11484C (.ZN(g11484C),.A2(g11461C),.A1(g6639C));
OR2_X1 U_g5842C (.ZN(g5842C),.A2(g3979C),.A1(g5618C));
OR4_X1 U_I15200C (.ZN(I15200C),.A4(g9880C),.A3(g9848C),.A2(g9962C),.A1(g9837C));
OR2_X1 U_g11609C (.ZN(g11609C),.A2(g11559C),.A1(g11588C));
OR2_X1 U_g8940C (.ZN(g8940C),.A2(FE_OFN332_g8748C),.A1(g8793C));
OR2_X1 U_g11312C (.ZN(g11312C),.A2(g11101C),.A1(g11222C));
OR2_X1 U_g11608C (.ZN(g11608C),.A2(g11558C),.A1(g11587C));
OR2_X1 U_g6000C (.ZN(g6000C),.A2(g3912C),.A1(g5480C));
OR2_X1 U_g8428C (.ZN(g8428C),.A2(g8068C),.A1(g8382C));
OR2_X1 U_g8430C (.ZN(g8430C),.A2(g8070C),.A1(g8386C));
OR2_X1 U_g9922C (.ZN(g9922C),.A2(g9705C),.A1(g9864C));
OR2_X1 U_g8247C (.ZN(g8247C),.A2(g7704C),.A1(g8010C));
OR2_X1 U_g3438C (.ZN(g3438C),.A2(g2944C),.A1(g2939C));
OR4_X1 U_I5576C (.ZN(I5576C),.A4(g444C),.A3(g440C),.A2(g435C),.A1(g431C));
OR2_X1 U_g6924C (.ZN(g6924C),.A2(g4261C),.A1(g6362C));
OR2_X1 U_g5405C (.ZN(g5405C),.A2(FE_OFN221_g3440C),.A1(g4476C));
OR2_X1 U_g8638C (.ZN(g8638C),.A2(g8461C),.A1(g8108C));
OR2_X1 U_g8609C (.ZN(g8609C),.A2(g8555C),.A1(g8408C));
OR2_X1 U_g9995C (.ZN(g9995C),.A2(I15200C),.A1(I15199C));
OR2_X1 U_g8883C (.ZN(g8883C),.A2(FE_OFN329_g8763C),.A1(g8838C));
OR4_X1 U_I15214C (.ZN(I15214C),.A4(g9831C),.A3(g9935C),.A2(g9906C),.A1(g8170C));
OR3_X1 U_g2538C (.ZN(g2538C),.A3(I5649C),.A2(g1458C),.A1(g1466C));
OR2_X1 U_g11329C (.ZN(g11329C),.A2(g11169C),.A1(g11302C));
OR2_X1 U_g4255C (.ZN(g4255C),.A2(g4047C),.A1(g4009C));
OR2_X1 U_g11328C (.ZN(g11328C),.A2(g11168C),.A1(g11299C));
OR3_X1 U_g9704C (.ZN(g9704C),.A3(I14835C),.A2(g9605C),.A1(g9385C));
OR4_X1 U_I5352C (.ZN(I5352C),.A4(g1117C),.A3(g1121C),.A2(g1125C),.A1(g1129C));
OR2_X1 U_g8774C (.ZN(g8774C),.A2(g8654C),.A1(g5499C));
OR3_X1 U_g9954C (.ZN(g9954C),.A3(g9803C),.A2(g9940C),.A1(g9946C));
OR2_X1 U_g10405C (.ZN(g10405C),.A2(g9291C),.A1(g10297C));
OR2_X1 U_g9363C (.ZN(g9363C),.A2(g9192C),.A1(g9205C));
OR2_X1 U_g5849C (.ZN(g5849C),.A2(g4144C),.A1(g4949C));
OR4_X1 U_I5599C (.ZN(I5599C),.A4(g501C),.A3(g506C),.A2(g511C),.A1(g516C));
OR2_X1 U_g7204C (.ZN(g7204C),.A2(I9717C),.A1(g6645C));
OR2_X1 U_g7300C (.ZN(g7300C),.A2(g6326C),.A1(g7139C));
OR2_X1 U_g4293C (.ZN(g4293C),.A2(g4068C),.A1(g4064C));
OR2_X1 U_g9912C (.ZN(g9912C),.A2(g9690C),.A1(g9847C));
OR2_X1 U_g6533C (.ZN(g6533C),.A2(g5002C),.A1(g5771C));
OR2_X1 U_g8816C (.ZN(g8816C),.A2(g8731C),.A1(g7951C));
OR2_X1 U_g9929C (.ZN(g9929C),.A2(g9718C),.A1(g9871C));
OR2_X1 U_g5819C (.ZN(g5819C),.A2(g4876C),.A1(g5625C));
OR3_X1 U_I14831C (.ZN(I14831C),.A3(g9586C),.A2(g9622C),.A1(g9613C));
OR2_X1 U_g5852C (.ZN(g5852C),.A2(g3989C),.A1(g5632C));
OR2_X1 U_g8263C (.ZN(g8263C),.A2(g7720C),.A1(g8032C));
OR2_X1 U_g3431C (.ZN(g3431C),.A2(g2957C),.A1(g2951C));
OR2_X1 U_g8631C (.ZN(g8631C),.A2(g7449C),.A1(g8474C));
OR2_X1 U_g6922C (.ZN(g6922C),.A2(g5694C),.A1(g6352C));
OR2_X1 U_g8817C (.ZN(g8817C),.A2(g8732C),.A1(g7954C));
OR4_X1 U_g9735C (.ZN(g9735C),.A4(g9387C),.A3(g9384C),.A2(g9651C),.A1(g9649C));
OR2_X1 U_g8605C (.ZN(g8605C),.A2(g8553C),.A1(g8404C));
OR2_X1 U_g11263C (.ZN(g11263C),.A2(g11025C),.A1(g11187C));
OR2_X1 U_g6739C (.ZN(g6739C),.A2(g5780C),.A1(g5769C));
OR2_X1 U_g11332C (.ZN(g11332C),.A2(g11172C),.A1(g11273C));
OR2_X1 U_g7143C (.ZN(g7143C),.A2(I9717C),.A1(g6619C));
OR2_X1 U_g6479C (.ZN(g6479C),.A2(g4968C),.A1(g5707C));
OR4_X1 U_I15048C (.ZN(I15048C),.A4(FE_OFN35_g9785C),.A3(FE_OFN61_g9624C),.A2(g9680C),.A1(FE_OFN90_I11360C));
OR2_X1 U_g6501C (.ZN(g6501C),.A2(g4987C),.A1(g5726C));
OR3_X1 U_g9702C (.ZN(g9702C),.A3(I14831C),.A2(g9647C),.A1(g9365C));
OR2_X1 U_g11221C (.ZN(g11221C),.A2(g11007C),.A1(g11146C));
OR3_X1 U_g9952C (.ZN(g9952C),.A3(g9815C),.A2(g9938C),.A1(g9944C));
OR2_X1 U_g11613C (.ZN(g11613C),.A2(g11591C),.A1(g11600C));
OR2_X1 U_g7621C (.ZN(g7621C),.A2(g6994C),.A1(g5108C));
OR2_X1 U_g3399C (.ZN(g3399C),.A2(g2940C),.A1(g2918C));
OR2_X1 U_g11605C (.ZN(g11605C),.A2(g11555C),.A1(g11584C));
OR2_X1 U_g4274C (.ZN(g4274C),.A2(g4058C),.A1(g4054C));
OR3_X1 U_I14602C (.ZN(I14602C),.A3(g9192C),.A2(FE_OFN42_g9205C),.A1(g8995C));
OR4_X1 U_I15033C (.ZN(I15033C),.A4(FE_OFN35_g9785C),.A3(FE_OFN61_g9624C),.A2(FE_OFN33_g9454C),.A1(FE_OFN90_I11360C));
OR2_X1 U_g10717C (.ZN(g10717C),.A2(g10705C),.A1(g6235C));
OR3_X1 U_I5629C (.ZN(I5629C),.A3(g837C),.A2(g841C),.A1(g845C));
OR2_X1 U_g9925C (.ZN(g9925C),.A2(g9712C),.A1(g9867C));
OR2_X1 U_g3819C (.ZN(g3819C),.A2(g9C),.A1(g3275C));
OR2_X1 U_g6912C (.ZN(g6912C),.A2(g4235C),.A1(g6350C));
OR2_X1 U_g10723C (.ZN(g10723C),.A2(g10633C),.A1(g4952C));
OR2_X1 U_g6929C (.ZN(g6929C),.A2(g5704C),.A1(g6360C));
OR2_X1 U_g10646C (.ZN(g10646C),.A2(g7739C),.A1(g10625C));
OR2_X1 U_g9516C (.ZN(g9516C),.A2(FE_OFN44_g9125C),.A1(FE_OFN47_g9151C));
OR2_X1 U_g6626C (.ZN(g6626C),.A2(g123C),.A1(g5934C));
OR4_X1 U_I6350C (.ZN(I6350C),.A4(g2419C),.A3(g2433C),.A2(g2437C),.A1(g2445C));
OR2_X1 U_g11325C (.ZN(g11325C),.A2(g11165C),.A1(g11295C));
OR4_X1 U_I5366C (.ZN(I5366C),.A4(g1296C),.A3(g1292C),.A2(g1284C),.A1(g1280C));
OR3_X1 U_I5649C (.ZN(I5649C),.A3(g1482C),.A2(g1486C),.A1(g1499C));
OR2_X1 U_g6894C (.ZN(g6894C),.A2(g4868C),.A1(g6763C));
OR3_X1 U_g9738C (.ZN(g9738C),.A3(g9506C),.A2(g9447C),.A1(g9417C));
OR2_X1 U_g8383C (.ZN(g8383C),.A2(g5051C),.A1(g8163C));
OR2_X1 U_g8779C (.ZN(g8779C),.A2(g8663C),.A1(g5530C));
OR2_X1 U_g8161C (.ZN(g8161C),.A2(g7185C),.A1(g8005C));
OR2_X2 U_g8451C (.ZN(g8451C),.A2(g8366C),.A1(FE_OFN221_g3440C));
OR2_X1 U_g9915C (.ZN(g9915C),.A2(g9693C),.A1(g9853C));
OR4_X1 U_g2316C (.ZN(g2316C),.A4(I5366C),.A3(g1270C),.A2(g1304C),.A1(g1300C));
OR2_X1 U_g5576C (.ZN(g5576C),.A2(FE_OFN204_g3664C),.A1(g4675C));
OR2_X1 U_g10857C (.ZN(g10857C),.A2(g10738C),.A1(g6090C));
OR2_X1 U_g10793C (.ZN(g10793C),.A2(g10763C),.A1(g6194C));
OR2_X1 U_g7511C (.ZN(g7511C),.A2(g6438C),.A1(g6890C));
OR2_X1 U_g8944C (.ZN(g8944C),.A2(FE_OFN332_g8748C),.A1(g8799C));
OR2_X1 U_g10765C (.ZN(g10765C),.A2(g10680C),.A1(g5492C));
OR2_X1 U_g10549C (.ZN(g10549C),.A2(g10451C),.A1(g4271C));
OR2_X1 U_g7092C (.ZN(g7092C),.A2(g5902C),.A1(g6540C));
OR2_X1 U_g11604C (.ZN(g11604C),.A2(g11554C),.A1(g11583C));
OR2_X1 U_g8434C (.ZN(g8434C),.A2(g8074C),.A1(g8400C));
OR2_X1 U_g6546C (.ZN(g6546C),.A2(g5026C),.A1(g5796C));
OR2_X1 U_g3354C (.ZN(g3354C),.A2(g1216C),.A1(g3121C));
OR2_X1 U_g9928C (.ZN(g9928C),.A2(g9717C),.A1(g9870C));
OR2_X1 U_g11262C (.ZN(g11262C),.A2(g11024C),.A1(g11240C));
OR4_X1 U_g9785C (.ZN(g9785C),.A4(g9363C),.A3(g9388C),.A2(g8995C),.A1(g9010C));
OR2_X1 U_g5867C (.ZN(g5867C),.A2(g4921C),.A1(FE_OFN221_g3440C));
OR2_X1 U_g8210C (.ZN(g8210C),.A2(g7692C),.A1(g7466C));
OR2_X1 U_g10533C (.ZN(g10533C),.A2(g10449C),.A1(g4437C));
OR2_X1 U_g9563C (.ZN(g9563C),.A2(g9030C),.A1(FE_OFN56_g9052C));
OR2_X1 U_g6906C (.ZN(g6906C),.A2(g5674C),.A1(g6791C));
OR2_X1 U_g7375C (.ZN(g7375C),.A2(g6745C),.A1(g7230C));
OR2_X1 U_g7651C (.ZN(g7651C),.A2(FE_OFN350_g3121C),.A1(g7135C));
OR4_X1 U_I5570C (.ZN(I5570C),.A4(g401C),.A3(g406C),.A2(g411C),.A1(g416C));
OR3_X1 U_g9731C (.ZN(g9731C),.A3(g9387C),.A2(g9364C),.A1(g9641C));
OR2_X1 U_g11247C (.ZN(g11247C),.A2(g10949C),.A1(g11097C));
OR4_X1 U_I15045C (.ZN(I15045C),.A4(FE_OFN35_g9785C),.A3(FE_OFN61_g9624C),.A2(g9676C),.A1(FE_OFN90_I11360C));
OR2_X1 U_g10856C (.ZN(g10856C),.A2(g10737C),.A1(g6083C));
OR2_X1 U_g7184C (.ZN(g7184C),.A2(g6047C),.A1(g6625C));
OR2_X1 U_g11612C (.ZN(g11612C),.A2(g11590C),.A1(g11599C));
OR2_X1 U_g7384C (.ZN(g7384C),.A2(g6618C),.A1(g7088C));
OR2_X1 U_g11324C (.ZN(g11324C),.A2(g11164C),.A1(g11271C));
OR2_X1 U_g8922C (.ZN(g8922C),.A2(FE_OFN329_g8763C),.A1(g8822C));
OR4_X1 U_I5358C (.ZN(I5358C),.A4(g1275C),.A3(g1235C),.A2(g1240C),.A1(g1245C));
OR3_X1 U_g9955C (.ZN(g9955C),.A3(g9803C),.A2(g9941C),.A1(g9947C));
OR4_X1 U_g2501C (.ZN(g2501C),.A4(I5576C),.A3(g421C),.A2(g452C),.A1(g448C));
OR2_X1 U_g7231C (.ZN(g7231C),.A2(g6087C),.A1(g6673C));
OR2_X1 U_g6078C (.ZN(g6078C),.A2(g5256C),.A1(g4503C));
OR2_X1 U_g6478C (.ZN(g6478C),.A2(g4967C),.A1(g5706C));
OR2_X1 U_g6907C (.ZN(g6907C),.A2(g5675C),.A1(g6792C));
OR2_X1 U_g6035C (.ZN(g6035C),.A2(g3974C),.A1(g5518C));
OR2_X1 U_g8937C (.ZN(g8937C),.A2(FE_OFN332_g8748C),.A1(g8786C));
OR2_X1 U_g7742C (.ZN(g7742C),.A2(g6743C),.A1(g7217C));
OR2_X1 U_g10722C (.ZN(g10722C),.A2(g10671C),.A1(g10308C));
OR2_X1 U_g9918C (.ZN(g9918C),.A2(g9698C),.A1(g9858C));
OR2_X1 U_g5403C (.ZN(g5403C),.A2(g3695C),.A1(g4486C));
OR2_X1 U_g7926C (.ZN(g7926C),.A2(g6892C),.A1(g7435C));
OR2_X1 U_g6915C (.ZN(g6915C),.A2(g5686C),.A1(g6347C));
OR2_X1 U_g5841C (.ZN(g5841C),.A2(g4230C),.A1(g4914C));
OR4_X1 U_I15220C (.ZN(I15220C),.A4(g9877C),.A3(g9857C),.A2(g9966C),.A1(g9841C));
OR2_X1 U_g10529C (.ZN(g10529C),.A2(I16161C),.A1(I16160C));
OR2_X1 U_g11246C (.ZN(g11246C),.A2(g10948C),.A1(g11094C));
OR2_X1 U_g6002C (.ZN(g6002C),.A2(g4827C),.A1(g5489C));
OR2_X1 U_g7712C (.ZN(g7712C),.A2(FE_OFN350_g3121C),.A1(g7125C));
OR2_X1 U_g8810C (.ZN(g8810C),.A2(g8720C),.A1(g7933C));
OR2_X1 U_g9921C (.ZN(g9921C),.A2(g9703C),.A1(g9862C));
OR2_X1 U_g8432C (.ZN(g8432C),.A2(g8072C),.A1(g8389C));
OR4_X1 U_I15172C (.ZN(I15172C),.A4(g9874C),.A3(g9861C),.A2(g9959C),.A1(g9843C));
OR3_X1 U_I14822C (.ZN(I14822C),.A3(g9582C),.A2(g9604C),.A1(g9597C));
OR2_X1 U_g6928C (.ZN(g6928C),.A2(g5703C),.A1(g6359C));
OR2_X1 U_g8157C (.ZN(g8157C),.A2(g7623C),.A1(FE_OFN192_g6488C));
OR2_X1 U_g6930C (.ZN(g6930C),.A2(g4269C),.A1(g6364C));
OR2_X1 U_g7660C (.ZN(g7660C),.A2(g5867C),.A1(g7059C));
OR2_X1 U_g6899C (.ZN(g6899C),.A2(g32C),.A1(g6463C));
OR2_X1 U_g9392C (.ZN(g9392C),.A2(g9324C),.A1(g9328C));
OR2_X1 U_g11318C (.ZN(g11318C),.A2(g11104C),.A1(g11228C));
OR3_X1 U_I16427C (.ZN(I16427C),.A3(g10382C),.A2(g10383C),.A1(g10683C));
OR2_X1 U_g11227C (.ZN(g11227C),.A2(g11010C),.A1(g11151C));
OR2_X1 U_g11058C (.ZN(g11058C),.A2(g5280C),.A1(g10933C));
OR4_X1 U_I5351C (.ZN(I5351C),.A4(g1133C),.A3(g1137C),.A2(g1141C),.A1(g1145C));
OR3_X1 U_g9708C (.ZN(g9708C),.A3(g9646C),.A2(g9389C),.A1(g9653C));
OR2_X1 U_g6071C (.ZN(g6071C),.A2(g4505C),.A1(g5228C));
OR2_X1 U_g9911C (.ZN(g9911C),.A2(g9689C),.A1(g9846C));
OR2_X1 U_g7102C (.ZN(g7102C),.A2(g5915C),.A1(g6550C));
OR2_X1 U_g7302C (.ZN(g7302C),.A2(g6328C),.A1(g7141C));
OR2_X1 U_g6038C (.ZN(g6038C),.A2(g3979C),.A1(g5528C));
OR2_X1 U_g4239C (.ZN(g4239C),.A2(g4008C),.A1(g4000C));
OR2_X1 U_g8646C (.ZN(g8646C),.A2(g8547C),.A1(g8224C));
OR2_X1 U_g9974C (.ZN(g9974C),.A2(I15177C),.A1(I15176C));
OR2_X1 U_g5823C (.ZN(g5823C),.A2(g4882C),.A1(g5631C));
OR2_X1 U_g6918C (.ZN(g6918C),.A2(g4252C),.A1(g6358C));
OR2_X1 U_g7265C (.ZN(g7265C),.A2(g6204C),.A1(g6756C));
OR4_X1 U_I5804C (.ZN(I5804C),.A4(g2104C),.A3(g2106C),.A2(g2109C),.A1(g2111C));
OR2_X1 U_g5851C (.ZN(g5851C),.A2(g4253C),.A1(g4941C));
OR2_X1 U_g11481C (.ZN(g11481C),.A2(g11458C),.A1(g6624C));
OR2_X1 U_g10336C (.ZN(g10336C),.A2(g9097C),.A1(g10230C));
OR2_X1 U_g7296C (.ZN(g7296C),.A2(g6322C),.A1(g7131C));
OR2_X1 U_g4300C (.ZN(g4300C),.A2(g1212C),.A1(g3546C));
OR2_X1 U_g8647C (.ZN(g8647C),.A2(g8470C),.A1(g8130C));
NAND2_X1 U_g8546C (.ZN(g8546C),.A2(g8390C),.A1(g3983C));
NAND2_X1 U_g2516C (.ZN(g2516C),.A2(I5613C),.A1(I5612C));
NAND2_X1 U_g2987C (.ZN(g2987C),.A2(g883C),.A1(g2481C));
NAND2_X1 U_I5593C (.ZN(I5593C),.A2(I5591C),.A1(g1703C));
NAND2_X1 U_g8970C (.ZN(g8970C),.A2(g8839C),.A1(g5548C));
NAND2_X1 U_I10519C (.ZN(I10519C),.A2(g822C),.A1(g6231C));
NAND2_X1 U_I11279C (.ZN(I11279C),.A2(I11278C),.A1(g305C));
NAND4_X1 U_g7990C (.ZN(g7990C),.A4(g7550C),.A3(g7562C),.A2(FE_OFN80_g2175C),.A1(FE_OFN88_g2178C));
NAND2_X1 U_I11278C (.ZN(I11278C),.A2(g6485C),.A1(g305C));
NAND2_X1 U_g3978C (.ZN(g3978C),.A2(g1822C),.A1(g3207C));
NAND2_X1 U_I5264C (.ZN(I5264C),.A2(I5263C),.A1(g456C));
NAND2_X1 U_I8640C (.ZN(I8640C),.A2(g516C),.A1(g4278C));
NAND2_X1 U_I6761C (.ZN(I6761C),.A2(I6760C),.A1(g2943C));
NAND2_X1 U_I17400C (.ZN(I17400C),.A2(g11416C),.A1(g11418C));
NAND2_X1 U_I5450C (.ZN(I5450C),.A2(I5449C),.A1(g1235C));
NAND2_X1 U_I16060C (.ZN(I16060C),.A2(I16058C),.A1(g10441C));
NAND2_X1 U_I6746C (.ZN(I6746C),.A2(g1453C),.A1(g2938C));
NAND2_X1 U_I11975C (.ZN(I11975C),.A2(I11973C),.A1(g1462C));
NAND2_X1 U_I12136C (.ZN(I12136C),.A2(g131C),.A1(g6038C));
NAND2_X1 U_I11937C (.ZN(I11937C),.A2(I11935C),.A1(g1458C));
NAND2_X1 U_g2959C (.ZN(g2959C),.A2(I6168C),.A1(I6167C));
NAND2_X1 U_I5878C (.ZN(I5878C),.A2(g2115C),.A1(g2120C));
NAND2_X1 U_g2517C (.ZN(g2517C),.A2(I5620C),.A1(I5619C));
NAND2_X1 U_g5552C (.ZN(g5552C),.A2(FE_OFN223_g4401C),.A1(g4777C));
NAND2_X1 U_I6468C (.ZN(I6468C),.A2(I6467C),.A1(g23C));
NAND2_X1 U_I8796C (.ZN(I8796C),.A2(I8795C),.A1(g4672C));
NAND2_X1 U_g10392C (.ZN(g10392C),.A2(I15892C),.A1(I15891C));
NAND2_X1 U_I5611C (.ZN(I5611C),.A2(g1284C),.A1(g1280C));
NAND2_X1 U_g8738C (.ZN(g8738C),.A2(FE_OFN200_g4921C),.A1(g8688C));
NAND2_X1 U_I6716C (.ZN(I6716C),.A2(I6714C),.A1(g201C));
NAND2_X1 U_g2310C (.ZN(g2310C),.A2(g605C),.A1(g591C));
NAND2_X1 U_I7685C (.ZN(I7685C),.A2(I7683C),.A1(g3460C));
NAND2_X1 U_g3056C (.ZN(g3056C),.A2(g599C),.A1(g2374C));
NAND2_X1 U_I12108C (.ZN(I12108C),.A2(I12106C),.A1(g135C));
NAND3_X1 U_g3529C (.ZN(g3529C),.A3(g2325C),.A2(g3062C),.A1(g2310C));
NAND2_X1 U_I6747C (.ZN(I6747C),.A2(I6746C),.A1(g2938C));
NAND2_X1 U_g2236C (.ZN(g2236C),.A2(I5231C),.A1(I5230C));
NAND2_X1 U_g7584C (.ZN(g7584C),.A2(I12076C),.A1(I12075C));
NAND2_X1 U_I15870C (.ZN(I15870C),.A2(FE_OFN239_g1796C),.A1(g10291C));
NAND2_X1 U_I16067C (.ZN(I16067C),.A2(I16065C),.A1(FE_OFN237_g1806C));
NAND2_X1 U_I7562C (.ZN(I7562C),.A2(g654C),.A1(g3533C));
NAND2_X1 U_I13531C (.ZN(I13531C),.A2(I13529C),.A1(g8253C));
NAND2_X1 U_I8797C (.ZN(I8797C),.A2(I8795C),.A1(g1145C));
NAND2_X1 U_I17584C (.ZN(I17584C),.A2(g11515C),.A1(g11217C));
NAND2_X1 U_I11936C (.ZN(I11936C),.A2(I11935C),.A1(g5857C));
NAND2_X1 U_I15257C (.ZN(I15257C),.A2(I15256C),.A1(g9974C));
NAND2_X1 U_g8402C (.ZN(g8402C),.A2(I13506C),.A1(I13505C));
NAND3_X1 U_g8824C (.ZN(g8824C),.A3(g8512C),.A2(g8501C),.A1(g8502C));
NAND2_X1 U_I6186C (.ZN(I6186C),.A2(g466C),.A1(g2511C));
NAND2_X1 U_g11496C (.ZN(g11496C),.A2(I17505C),.A1(I17504C));
NAND2_X1 U_I16001C (.ZN(I16001C),.A2(I15999C),.A1(FE_OFN247_g1771C));
NAND2_X1 U_I6125C (.ZN(I6125C),.A2(I6124C),.A1(g2215C));
NAND2_X1 U_I11909C (.ZN(I11909C),.A2(I11907C),.A1(g1474C));
NAND2_X1 U_I12040C (.ZN(I12040C),.A2(I12038C),.A1(g1466C));
NAND2_X1 U_I13909C (.ZN(I13909C),.A2(I13907C),.A1(g1432C));
NAND2_X1 U_g3625C (.ZN(g3625C),.A2(I6772C),.A1(I6771C));
NAND2_X1 U_I11908C (.ZN(I11908C),.A2(I11907C),.A1(g5838C));
NAND2_X1 U_g10470C (.ZN(g10470C),.A2(I16009C),.A1(I16008C));
NAND2_X1 U_I13908C (.ZN(I13908C),.A2(I13907C),.A1(g8265C));
NAND2_X1 U_g3813C (.ZN(g3813C),.A2(I7035C),.A1(I7034C));
NAND2_X1 U_I8650C (.ZN(I8650C),.A2(g778C),.A1(g4824C));
NAND2_X1 U_g6207C (.ZN(g6207C),.A2(I9948C),.A1(I9947C));
NAND2_X1 U_I16066C (.ZN(I16066C),.A2(I16065C),.A1(g10428C));
NAND2_X1 U_g2948C (.ZN(g2948C),.A2(I6145C),.A1(I6144C));
NAND2_X1 U_I11242C (.ZN(I11242C),.A2(I11241C),.A1(g6760C));
NAND2_X1 U_g10467C (.ZN(g10467C),.A2(I15994C),.A1(I15993C));
NAND2_X1 U_I6187C (.ZN(I6187C),.A2(I6186C),.A1(g2511C));
NAND2_X1 U_g6488C (.ZN(g6488C),.A2(g6019C),.A1(g6027C));
NAND2_X1 U_I5500C (.ZN(I5500C),.A2(g1007C),.A1(g1255C));
NAND2_X1 U_I11974C (.ZN(I11974C),.A2(I11973C),.A1(g5852C));
NAND2_X1 U_I12062C (.ZN(I12062C),.A2(I12060C),.A1(g1478C));
NAND2_X1 U_g5300C (.ZN(g5300C),.A2(I8772C),.A1(I8771C));
NAND2_X1 U_I5184C (.ZN(I5184C),.A2(g1515C),.A1(g1415C));
NAND2_X1 U_I13293C (.ZN(I13293C),.A2(g8161C),.A1(g1882C));
NAND2_X1 U_I6200C (.ZN(I6200C),.A2(I6199C),.A1(g2525C));
NAND2_X1 U_I13265C (.ZN(I13265C),.A2(g8154C),.A1(g1909C));
NAND2_X1 U_I5024C (.ZN(I5024C),.A2(I5023C),.A1(g995C));
NAND2_X1 U_I7863C (.ZN(I7863C),.A2(g774C),.A1(g4099C));
NAND2_X1 U_g8705C (.ZN(g8705C),.A2(I13992C),.A1(I13991C));
NAND2_X1 U_g8471C (.ZN(g8471C),.A2(I13661C),.A1(I13660C));
NAND2_X1 U_I15256C (.ZN(I15256C),.A2(g9968C),.A1(g9974C));
NAND2_X1 U_I6145C (.ZN(I6145C),.A2(I6143C),.A1(g646C));
NAND2_X1 U_I13992C (.ZN(I13992C),.A2(I13990C),.A1(g8688C));
NAND2_X1 U_I11510C (.ZN(I11510C),.A2(I11508C),.A1(FE_OFN237_g1806C));
NAND2_X1 U_g10853C (.ZN(g10853C),.A2(g5034C),.A1(g10731C));
NAND2_X1 U_I5231C (.ZN(I5231C),.A2(I5229C),.A1(g148C));
NAND2_X1 U_I12047C (.ZN(I12047C),.A2(I12045C),.A1(g1486C));
NAND2_X1 U_I10771C (.ZN(I10771C),.A2(I10769C),.A1(g1801C));
NAND2_X1 U_g10477C (.ZN(g10477C),.A2(I16046C),.A1(I16045C));
NAND2_X1 U_g7582C (.ZN(g7582C),.A2(I12062C),.A1(I12061C));
NAND2_X1 U_I5104C (.ZN(I5104C),.A2(g435C),.A1(g431C));
NAND2_X1 U_g8409C (.ZN(g8409C),.A2(I13531C),.A1(I13530C));
NAND2_X1 U_I6447C (.ZN(I6447C),.A2(FE_OFN236_g1776C),.A1(g2264C));
NAND2_X1 U_I4956C (.ZN(I4956C),.A2(I4954C),.A1(g327C));
NAND2_X1 U_I5613C (.ZN(I5613C),.A2(I5611C),.A1(g1284C));
NAND2_X1 U_I8481C (.ZN(I8481C),.A2(I8479C),.A1(g3530C));
NAND2_X1 U_g5278C (.ZN(g5278C),.A2(I8740C),.A1(I8739C));
NAND2_X1 U_I6880C (.ZN(I6880C),.A2(I6879C),.A1(g3301C));
NAND2_X1 U_I15431C (.ZN(I15431C),.A2(I15430C),.A1(g10001C));
NAND2_X1 U_g5548C (.ZN(g5548C),.A2(FE_OFN223_g4401C),.A1(g1840C));
NAND4_X1 U_g7671C (.ZN(g7671C),.A4(FE_OFN96_g2169C),.A3(FE_OFN91_g2172C),.A2(g2175C),.A1(g2178C));
NAND2_X1 U_I12020C (.ZN(I12020C),.A2(I12019C),.A1(g6049C));
NAND2_X1 U_g10665C (.ZN(g10665C),.A2(I16332C),.A1(I16331C));
NAND2_X1 U_I16469C (.ZN(I16469C),.A2(I16467C),.A1(g10518C));
NAND2_X1 U_I5014C (.ZN(I5014C),.A2(I5013C),.A1(g1007C));
NAND2_X1 U_I13523C (.ZN(I13523C),.A2(I13521C),.A1(g8249C));
NAND2_X1 U_I16039C (.ZN(I16039C),.A2(I16037C),.A1(FE_OFN252_g1791C));
NAND2_X1 U_I16468C (.ZN(I16468C),.A2(I16467C),.A1(g10716C));
NAND2_X1 U_I12046C (.ZN(I12046C),.A2(I12045C),.A1(g5814C));
NAND2_X1 U_g4476C (.ZN(g4476C),.A2(g3071C),.A1(g3807C));
NAND2_X1 U_g10476C (.ZN(g10476C),.A2(I16039C),.A1(I16038C));
NAND2_X1 U_I16038C (.ZN(I16038C),.A2(I16037C),.A1(g10363C));
NAND2_X1 U_I8676C (.ZN(I8676C),.A2(g1027C),.A1(g4374C));
NAND2_X1 U_I12113C (.ZN(I12113C),.A2(g162C),.A1(g6002C));
NAND2_X1 U_I8761C (.ZN(I8761C),.A2(g1129C),.A1(g4616C));
NAND2_X1 U_g3204C (.ZN(g3204C),.A2(g2061C),.A1(g2571C));
NAND2_X1 U_I15993C (.ZN(I15993C),.A2(I15992C),.A1(g10430C));
NAND2_X1 U_I5036C (.ZN(I5036C),.A2(I5034C),.A1(g1019C));
NAND2_X1 U_I14263C (.ZN(I14263C),.A2(g1814C),.A1(g8843C));
NAND2_X1 U_g8298C (.ZN(g8298C),.A2(I13250C),.A1(I13249C));
NAND2_X1 U_I5135C (.ZN(I5135C),.A2(g525C),.A1(g521C));
NAND2_X1 U_g2405C (.ZN(g2405C),.A2(I5486C),.A1(I5485C));
NAND2_X1 U_I7034C (.ZN(I7034C),.A2(I7033C),.A1(g3089C));
NAND2_X1 U_I15443C (.ZN(I15443C),.A2(I15441C),.A1(g10007C));
NAND2_X1 U_I6166C (.ZN(I6166C),.A2(g153C),.A1(g2236C));
NAND2_X1 U_I8624C (.ZN(I8624C),.A2(g511C),.A1(g4267C));
NAND2_X1 U_I16015C (.ZN(I16015C),.A2(g1781C),.A1(g10441C));
NAND2_X1 U_I8677C (.ZN(I8677C),.A2(I8676C),.A1(g4374C));
NAND2_X1 U_I8576C (.ZN(I8576C),.A2(I8575C),.A1(g4234C));
NAND2_X1 U_I14613C (.ZN(I14613C),.A2(I14612C),.A1(g9204C));
NAND2_X1 U_I8716C (.ZN(I8716C),.A2(I8715C),.A1(g4601C));
NAND2_X1 U_g3530C (.ZN(g3530C),.A2(I6716C),.A1(I6715C));
NAND2_X1 U_g8405C (.ZN(g8405C),.A2(I13515C),.A1(I13514C));
NAND4_X1 U_g4104C (.ZN(g4104C),.A4(g3200C),.A3(g2439C),.A2(g3247C),.A1(g3215C));
NAND2_X1 U_I12003C (.ZN(I12003C),.A2(I12002C),.A1(g5996C));
NAND2_X1 U_g2177C (.ZN(g2177C),.A2(I5128C),.A1(I5127C));
NAND2_X1 U_g3010C (.ZN(g3010C),.A2(g2399C),.A1(g2382C));
NAND2_X1 U_g5179C (.ZN(g5179C),.A2(I8577C),.A1(I8576C));
NAND2_X1 U_I17395C (.ZN(I17395C),.A2(I17393C),.A1(g11414C));
NAND2_X1 U_g7067C (.ZN(g7067C),.A2(I11280C),.A1(I11279C));
NAND4_X1 U_g7994C (.ZN(g7994C),.A4(g7550C),.A3(FE_OFN91_g2172C),.A2(g7574C),.A1(FE_OFN88_g2178C));
NAND2_X1 U_I6167C (.ZN(I6167C),.A2(I6166C),.A1(g2236C));
NAND2_X1 U_I5265C (.ZN(I5265C),.A2(I5263C),.A1(g461C));
NAND2_X1 U_I6989C (.ZN(I6989C),.A2(I6988C),.A1(g2760C));
NAND2_X1 U_I13274C (.ZN(I13274C),.A2(I13272C),.A1(g8158C));
NAND2_X1 U_I10507C (.ZN(I10507C),.A2(g786C),.A1(g6221C));
NAND2_X1 U_I13530C (.ZN(I13530C),.A2(I13529C),.A1(g704C));
NAND2_X1 U_I5164C (.ZN(I5164C),.A2(g1499C),.A1(g1508C));
NAND2_X1 U_g9107C (.ZN(g9107C),.A2(I14444C),.A1(I14443C));
NAND2_X1 U_I9559C (.ZN(I9559C),.A2(I9557C),.A1(g782C));
NAND2_X1 U_I8577C (.ZN(I8577C),.A2(I8575C),.A1(g496C));
NAND2_X1 U_g2510C (.ZN(g2510C),.A2(I5593C),.A1(I5592C));
NAND2_X1 U_g8177C (.ZN(g8177C),.A2(I13078C),.A1(I13077C));
NAND2_X1 U_I8717C (.ZN(I8717C),.A2(I8715C),.A1(g4052C));
NAND2_X1 U_I5296C (.ZN(I5296C),.A2(I5295C),.A1(g794C));
NAND2_X1 U_g5209C (.ZN(g5209C),.A2(I8626C),.A1(I8625C));
NAND4_X1 U_g7950C (.ZN(g7950C),.A4(FE_OFN96_g2169C),.A3(g7562C),.A2(g7574C),.A1(g6941C));
NAND2_X1 U_g2088C (.ZN(g2088C),.A2(I4912C),.A1(I4911C));
NAND2_X1 U_I16000C (.ZN(I16000C),.A2(I15999C),.A1(g10432C));
NAND2_X1 U_I5371C (.ZN(I5371C),.A2(g976C),.A1(g971C));
NAND2_X1 U_g2215C (.ZN(g2215C),.A2(I5186C),.A1(I5185C));
NAND2_X1 U_g7101C (.ZN(g7101C),.A2(g2364C),.A1(g6617C));
NAND2_X1 U_I5675C (.ZN(I5675C),.A2(g1223C),.A1(g1218C));
NAND2_X1 U_I8544C (.ZN(I8544C),.A2(I8543C),.A1(g4218C));
NAND2_X1 U_g6577C (.ZN(g6577C),.A2(I10521C),.A1(I10520C));
NAND2_X1 U_I5297C (.ZN(I5297C),.A2(I5295C),.A1(g798C));
NAND2_X1 U_I13537C (.ZN(I13537C),.A2(g8157C),.A1(g658C));
NAND2_X1 U_I13283C (.ZN(I13283C),.A2(g8159C),.A1(g1927C));
NAND2_X1 U_g4749C (.ZN(g4749C),.A2(g2061C),.A1(g3710C));
NAND2_X1 U_I11982C (.ZN(I11982C),.A2(I11980C),.A1(g1482C));
NAND2_X1 U_I8514C (.ZN(I8514C),.A2(I8513C),.A1(g4873C));
NAND2_X1 U_I13091C (.ZN(I13091C),.A2(I13089C),.A1(g1840C));
NAND2_X1 U_g2943C (.ZN(g2943C),.A2(I6126C),.A1(I6125C));
NAND2_X1 U_I15908C (.ZN(I15908C),.A2(I15906C),.A1(g10302C));
NAND2_X1 U_I6879C (.ZN(I6879C),.A2(g1351C),.A1(g3301C));
NAND2_X1 U_I8763C (.ZN(I8763C),.A2(I8761C),.A1(g1129C));
NAND2_X1 U_I5449C (.ZN(I5449C),.A2(g991C),.A1(g1235C));
NAND3_X1 U_g8825C (.ZN(g8825C),.A3(g8506C),.A2(g8738C),.A1(g8502C));
NAND2_X1 U_I16007C (.ZN(I16007C),.A2(FE_OFN236_g1776C),.A1(g10434C));
NAND2_X1 U_I5865C (.ZN(I5865C),.A2(g2105C),.A1(g2107C));
NAND2_X1 U_I5604C (.ZN(I5604C),.A2(g1153C),.A1(g1149C));
NAND2_X1 U_g2433C (.ZN(g2433C),.A2(I5518C),.A1(I5517C));
NAND2_X1 U_I6111C (.ZN(I6111C),.A2(I6109C),.A1(g1494C));
NAND2_X1 U_g2096C (.ZN(g2096C),.A2(I4930C),.A1(I4929C));
NAND2_X1 U_I13522C (.ZN(I13522C),.A2(I13521C),.A1(g695C));
NAND2_X1 U_I10770C (.ZN(I10770C),.A2(I10769C),.A1(g5944C));
NAND2_X1 U_g6027C (.ZN(g6027C),.A2(FE_OFN200_g4921C),.A1(g4566C));
NAND4_X1 U_g7992C (.ZN(g7992C),.A4(FE_OFN96_g2169C),.A3(FE_OFN91_g2172C),.A2(g7574C),.A1(FE_OFN88_g2178C));
NAND2_X1 U_I5539C (.ZN(I5539C),.A2(I5538C),.A1(g1270C));
NAND2_X1 U_I17394C (.ZN(I17394C),.A2(I17393C),.A1(g11415C));
NAND2_X1 U_I13553C (.ZN(I13553C),.A2(I13552C),.A1(g668C));
NAND2_X1 U_I8642C (.ZN(I8642C),.A2(I8640C),.A1(g516C));
NAND2_X1 U_g7573C (.ZN(g7573C),.A2(I12047C),.A1(I12046C));
NAND2_X1 U_g11416C (.ZN(g11416C),.A2(I17297C),.A1(I17296C));
NAND2_X1 U_g6003C (.ZN(g6003C),.A2(g5548C),.A1(g5552C));
NAND2_X1 U_g8934C (.ZN(g8934C),.A2(I14279C),.A1(I14278C));
NAND2_X1 U_I15992C (.ZN(I15992C),.A2(g2677C),.A1(g10430C));
NAND2_X1 U_I7683C (.ZN(I7683C),.A2(g3460C),.A1(g1023C));
NAND2_X1 U_I4910C (.ZN(I4910C),.A2(g318C),.A1(g386C));
NAND4_X1 U_g3209C (.ZN(g3209C),.A4(g2571C),.A3(g2564C),.A2(g2061C),.A1(g2550C));
NAND2_X1 U_I6794C (.ZN(I6794C),.A2(I6792C),.A1(g143C));
NAND2_X1 U_I10521C (.ZN(I10521C),.A2(I10519C),.A1(g822C));
NAND2_X1 U_I5486C (.ZN(I5486C),.A2(I5484C),.A1(g1011C));
NAND2_X1 U_I15442C (.ZN(I15442C),.A2(I15441C),.A1(g10013C));
NAND2_X1 U_g6858C (.ZN(g6858C),.A2(I10932C),.A1(I10931C));
NAND2_X1 U_I5185C (.ZN(I5185C),.A2(I5184C),.A1(g1415C));
NAND2_X1 U_g5304C (.ZN(g5304C),.A2(I8780C),.A1(I8779C));
NAND2_X1 U_g2354C (.ZN(g2354C),.A2(g1520C),.A1(g1515C));
NAND2_X1 U_I15615C (.ZN(I15615C),.A2(g10153C),.A1(g10043C));
NAND2_X1 U_I17281C (.ZN(I17281C),.A2(g11219C),.A1(g11221C));
NAND2_X1 U_I5470C (.ZN(I5470C),.A2(I5468C),.A1(g999C));
NAND2_X1 U_I11509C (.ZN(I11509C),.A2(I11508C),.A1(g6580C));
NAND2_X1 U_I5025C (.ZN(I5025C),.A2(I5023C),.A1(g1275C));
NAND2_X1 U_I11508C (.ZN(I11508C),.A2(g1806C),.A1(g6580C));
NAND2_X1 U_I15430C (.ZN(I15430C),.A2(g9995C),.A1(g10001C));
NAND2_X1 U_I14612C (.ZN(I14612C),.A2(g611C),.A1(g9204C));
NAND2_X1 U_g4675C (.ZN(g4675C),.A2(g3247C),.A1(g4073C));
NAND2_X1 U_I14272C (.ZN(I14272C),.A2(I14270C),.A1(g1822C));
NAND2_X1 U_g2979C (.ZN(g2979C),.A2(I6209C),.A1(I6208C));
NAND2_X1 U_I17290C (.ZN(I17290C),.A2(I17288C),.A1(g11223C));
NAND2_X1 U_g5269C (.ZN(g5269C),.A2(I8717C),.A1(I8716C));
NAND2_X1 U_g4297C (.ZN(g4297C),.A2(I7564C),.A1(I7563C));
NAND2_X1 U_I12002C (.ZN(I12002C),.A2(g153C),.A1(g5996C));
NAND2_X1 U_I5006C (.ZN(I5006C),.A2(I5005C),.A1(g421C));
NAND2_X1 U_I12128C (.ZN(I12128C),.A2(I12126C),.A1(g170C));
NAND2_X1 U_I5105C (.ZN(I5105C),.A2(I5104C),.A1(g431C));
NAND2_X1 U_I6323C (.ZN(I6323C),.A2(I6322C),.A1(g2050C));
NAND2_X1 U_g7588C (.ZN(g7588C),.A2(I12094C),.A1(I12093C));
NAND2_X1 U_I6666C (.ZN(I6666C),.A2(I6664C),.A1(g2776C));
NAND2_X1 U_g3623C (.ZN(g3623C),.A2(I6762C),.A1(I6761C));
NAND2_X1 U_I5373C (.ZN(I5373C),.A2(I5371C),.A1(g976C));
NAND2_X1 U_I8529C (.ZN(I8529C),.A2(I8527C),.A1(g481C));
NAND2_X1 U_I5283C (.ZN(I5283C),.A2(I5282C),.A1(g758C));
NAND2_X1 U_I7224C (.ZN(I7224C),.A2(I7223C),.A1(g2981C));
NAND2_X1 U_I5007C (.ZN(I5007C),.A2(I5005C),.A1(g312C));
NAND2_X1 U_I5459C (.ZN(I5459C),.A2(g1003C),.A1(g1240C));
NAND2_X1 U_I17297C (.ZN(I17297C),.A2(I17295C),.A1(g11227C));
NAND3_X1 U_g8746C (.ZN(g8746C),.A3(g46C),.A2(g47C),.A1(g8617C));
NAND2_X1 U_I6143C (.ZN(I6143C),.A2(g646C),.A1(g1976C));
NAND2_X1 U_I5015C (.ZN(I5015C),.A2(I5013C),.A1(g1011C));
NAND2_X1 U_g8932C (.ZN(g8932C),.A2(I14265C),.A1(I14264C));
NAND2_X1 U_I16073C (.ZN(I16073C),.A2(I16072C),.A1(g845C));
NAND2_X1 U_I6988C (.ZN(I6988C),.A2(g986C),.A1(g2760C));
NAND2_X1 U_g3205C (.ZN(g3205C),.A2(g2571C),.A1(g1814C));
NAND2_X1 U_I8652C (.ZN(I8652C),.A2(I8650C),.A1(g778C));
NAND2_X1 U_I9558C (.ZN(I9558C),.A2(I9557C),.A1(g5598C));
NAND2_X1 U_I5203C (.ZN(I5203C),.A2(I5202C),.A1(g369C));
NAND2_X1 U_g7533C (.ZN(g7533C),.A2(I11937C),.A1(I11936C));
NAND2_X1 U_g3634C (.ZN(g3634C),.A2(I6807C),.A1(I6806C));
NAND2_X1 U_I6792C (.ZN(I6792C),.A2(g143C),.A1(g2959C));
NAND2_X1 U_g3304C (.ZN(g3304C),.A2(I6469C),.A1(I6468C));
NAND2_X1 U_I12145C (.ZN(I12145C),.A2(I12143C),.A1(g158C));
NAND2_X1 U_g7596C (.ZN(g7596C),.A2(I12128C),.A1(I12127C));
NAND2_X1 U_I13302C (.ZN(I13302C),.A2(I13300C),.A1(g8162C));
NAND2_X1 U_I5502C (.ZN(I5502C),.A2(I5500C),.A1(g1007C));
NAND2_X1 U_I9574C (.ZN(I9574C),.A2(g818C),.A1(g5608C));
NAND2_X1 U_g3273C (.ZN(g3273C),.A2(I6449C),.A1(I6448C));
NAND2_X1 U_I8670C (.ZN(I8670C),.A2(I8669C),.A1(g4831C));
NAND2_X1 U_I7035C (.ZN(I7035C),.A2(I7033C),.A1(g1868C));
NAND2_X1 U_I15453C (.ZN(I15453C),.A2(I15451C),.A1(g10019C));
NAND2_X1 U_I8625C (.ZN(I8625C),.A2(I8624C),.A1(g4267C));
NAND2_X1 U_I7876C (.ZN(I7876C),.A2(I7875C),.A1(g4109C));
NAND2_X1 U_I14203C (.ZN(I14203C),.A2(I14202C),.A1(g8825C));
NAND2_X1 U_I15607C (.ZN(I15607C),.A2(g10144C),.A1(g10149C));
NAND2_X1 U_g2274C (.ZN(g2274C),.A2(I5325C),.A1(I5324C));
NAND2_X1 U_I8740C (.ZN(I8740C),.A2(I8738C),.A1(g1121C));
NAND2_X1 U_I17296C (.ZN(I17296C),.A2(I17295C),.A1(g11229C));
NAND2_X1 U_g10507C (.ZN(g10507C),.A2(g5859C),.A1(g10434C));
NAND2_X1 U_g2325C (.ZN(g2325C),.A2(g617C),.A1(g611C));
NAND2_X1 U_I8606C (.ZN(I8606C),.A2(I8604C),.A1(g506C));
NAND2_X1 U_I12087C (.ZN(I12087C),.A2(I12085C),.A1(g1470C));
NAND2_X1 U_I13249C (.ZN(I13249C),.A2(I13248C),.A1(g1891C));
NAND2_X1 U_I13248C (.ZN(I13248C),.A2(g8148C),.A1(g1891C));
NAND2_X1 U_I13552C (.ZN(I13552C),.A2(g8262C),.A1(g668C));
NAND2_X1 U_g2106C (.ZN(g2106C),.A2(I4980C),.A1(I4979C));
NAND2_X1 U_I12069C (.ZN(I12069C),.A2(I12067C),.A1(g139C));
NAND2_X1 U_g9204C (.ZN(g9204C),.A2(g8942C),.A1(g6019C));
NAND2_X1 U_I12068C (.ZN(I12068C),.A2(I12067C),.A1(g6045C));
NAND2_X1 U_I17503C (.ZN(I17503C),.A2(g5269C),.A1(g11430C));
NAND2_X1 U_I7877C (.ZN(I7877C),.A2(I7875C),.A1(g810C));
NAND2_X1 U_I5165C (.ZN(I5165C),.A2(I5164C),.A1(g1508C));
NAND2_X1 U_g6740C (.ZN(g6740C),.A2(g2550C),.A1(g6131C));
NAND2_X1 U_I6289C (.ZN(I6289C),.A2(I6287C),.A1(g981C));
NAND2_X1 U_I6777C (.ZN(I6777C),.A2(g650C),.A1(g2892C));
NAND2_X1 U_g5171C (.ZN(g5171C),.A2(I8563C),.A1(I8562C));
NAND2_X1 U_I15891C (.ZN(I15891C),.A2(I15890C),.A1(g853C));
NAND2_X1 U_I13090C (.ZN(I13090C),.A2(I13089C),.A1(g8006C));
NAND2_X1 U_g11474C (.ZN(g11474C),.A2(I17461C),.A1(I17460C));
NAND4_X1 U_g7942C (.ZN(g7942C),.A4(g7550C),.A3(g7562C),.A2(FE_OFN80_g2175C),.A1(g6941C));
NAND2_X1 U_I5538C (.ZN(I5538C),.A2(g1023C),.A1(g1270C));
NAND2_X1 U_I7563C (.ZN(I7563C),.A2(I7562C),.A1(g3533C));
NAND2_X1 U_I13513C (.ZN(I13513C),.A2(g8248C),.A1(g686C));
NAND2_X1 U_g2107C (.ZN(g2107C),.A2(I4987C),.A1(I4986C));
NAND2_X1 U_g2223C (.ZN(g2223C),.A2(I5204C),.A1(I5203C));
NAND2_X1 U_I13505C (.ZN(I13505C),.A2(I13504C),.A1(g677C));
NAND2_X1 U_I6209C (.ZN(I6209C),.A2(I6207C),.A1(g802C));
NAND2_X1 U_I12086C (.ZN(I12086C),.A2(I12085C),.A1(g5842C));
NAND2_X1 U_I8545C (.ZN(I8545C),.A2(I8543C),.A1(g486C));
NAND2_X1 U_I8180C (.ZN(I8180C),.A2(I8178C),.A1(FE_OFN253_g1786C));
NAND2_X1 U_g2115C (.ZN(g2115C),.A2(I5015C),.A1(I5014C));
NAND2_X1 U_I8591C (.ZN(I8591C),.A2(I8589C),.A1(g501C));
NAND2_X1 U_I10931C (.ZN(I10931C),.A2(I10930C),.A1(g5863C));
NAND2_X1 U_I17402C (.ZN(I17402C),.A2(I17400C),.A1(g11416C));
NAND2_X1 U_g8307C (.ZN(g8307C),.A2(I13295C),.A1(I13294C));
NAND2_X1 U_I12144C (.ZN(I12144C),.A2(I12143C),.A1(g6000C));
NAND2_X1 U_I10520C (.ZN(I10520C),.A2(I10519C),.A1(g6231C));
NAND2_X1 U_I5263C (.ZN(I5263C),.A2(FE_OFN254_g461C),.A1(g456C));
NAND2_X1 U_g8757C (.ZN(g8757C),.A2(FE_OFN223_g4401C),.A1(g8599C));
NAND2_X1 U_I6714C (.ZN(I6714C),.A2(g201C),.A1(g2961C));
NAND2_X1 U_I14211C (.ZN(I14211C),.A2(I14209C),.A1(g599C));
NAND2_X1 U_I8515C (.ZN(I8515C),.A2(I8513C),.A1(g3513C));
NAND2_X1 U_g2272C (.ZN(g2272C),.A2(I5317C),.A1(I5316C));
NAND2_X1 U_I9946C (.ZN(I9946C),.A2(g1796C),.A1(g5233C));
NAND2_X1 U_I8750C (.ZN(I8750C),.A2(g1125C),.A1(g4613C));
NAND2_X1 U_I5605C (.ZN(I5605C),.A2(I5604C),.A1(g1149C));
NAND2_X1 U_g8880C (.ZN(g8880C),.A2(I14204C),.A1(I14203C));
NAND2_X1 U_I16051C (.ZN(I16051C),.A2(g10434C),.A1(g837C));
NAND2_X1 U_I16072C (.ZN(I16072C),.A2(g10438C),.A1(g845C));
NAND2_X1 U_g10440C (.ZN(g10440C),.A2(g6037C),.A1(g10360C));
NAND2_X1 U_g8612C (.ZN(g8612C),.A2(I13859C),.A1(I13858C));
NAND2_X1 U_I15872C (.ZN(I15872C),.A2(I15870C),.A1(FE_OFN239_g1796C));
NAND2_X1 U_I8528C (.ZN(I8528C),.A2(I8527C),.A1(g4879C));
NAND2_X1 U_g8629C (.ZN(g8629C),.A2(I13902C),.A1(I13901C));
NAND4_X1 U_g8542C (.ZN(g8542C),.A4(g8390C),.A3(g1814C),.A2(g1828C),.A1(g2571C));
NAND2_X1 U_I9947C (.ZN(I9947C),.A2(I9946C),.A1(g5233C));
NAND2_X1 U_I6838C (.ZN(I6838C),.A2(I6836C),.A1(g806C));
NAND2_X1 U_g7583C (.ZN(g7583C),.A2(I12069C),.A1(I12068C));
NAND2_X1 U_g4803C (.ZN(g4803C),.A2(FE_OFN325_g18C),.A1(g3664C));
NAND2_X1 U_I17307C (.ZN(I17307C),.A2(I17305C),.A1(g11231C));
NAND2_X1 U_g4538C (.ZN(g4538C),.A2(g2399C),.A1(g3475C));
NAND2_X1 U_I15452C (.ZN(I15452C),.A2(I15451C),.A1(g10025C));
NAND2_X1 U_I13857C (.ZN(I13857C),.A2(g1448C),.A1(g8270C));
NAND2_X1 U_I14202C (.ZN(I14202C),.A2(g591C),.A1(g8825C));
NAND2_X1 U_I13765C (.ZN(I13765C),.A2(g8417C),.A1(g731C));
NAND2_X1 U_g2260C (.ZN(g2260C),.A2(I5297C),.A1(I5296C));
NAND4_X1 U_g7986C (.ZN(g7986C),.A4(g7550C),.A3(g2172C),.A2(FE_OFN80_g2175C),.A1(FE_OFN88_g2178C));
NAND2_X1 U_g5226C (.ZN(g5226C),.A2(I8671C),.A1(I8670C));
NAND2_X1 U_g8512C (.ZN(g8512C),.A2(g8366C),.A1(g3723C));
NAND2_X1 U_I16046C (.ZN(I16046C),.A2(I16044C),.A1(g10432C));
NAND2_X1 U_I13504C (.ZN(I13504C),.A2(g8247C),.A1(g677C));
NAND2_X1 U_g10447C (.ZN(g10447C),.A2(g5360C),.A1(g10363C));
NAND2_X1 U_g2167C (.ZN(g2167C),.A2(I5106C),.A1(I5105C));
NAND2_X1 U_I8804C (.ZN(I8804C),.A2(I8803C),.A1(g4677C));
NAND2_X1 U_g10472C (.ZN(g10472C),.A2(I16017C),.A1(I16016C));
NAND2_X1 U_I17487C (.ZN(I17487C),.A2(I17485C),.A1(g11474C));
NAND2_X1 U_I4995C (.ZN(I4995C),.A2(g309C),.A1(g416C));
NAND2_X1 U_I12093C (.ZN(I12093C),.A2(I12092C),.A1(g5810C));
NAND4_X1 U_g7987C (.ZN(g7987C),.A4(FE_OFN96_g2169C),.A3(g7562C),.A2(FE_OFN80_g2175C),.A1(FE_OFN88_g2178C));
NAND2_X1 U_g5227C (.ZN(g5227C),.A2(I8678C),.A1(I8677C));
NAND2_X1 U_I5126C (.ZN(I5126C),.A2(g1389C),.A1(g1386C));
NAND2_X1 U_g2321C (.ZN(g2321C),.A2(I5373C),.A1(I5372C));
NAND2_X1 U_g7547C (.ZN(g7547C),.A2(I11975C),.A1(I11974C));
NAND2_X1 U_I17306C (.ZN(I17306C),.A2(I17305C),.A1(g11232C));
NAND3_X1 U_g6548C (.ZN(g6548C),.A3(g6122C),.A2(g6124C),.A1(g826C));
NAND2_X1 U_I11995C (.ZN(I11995C),.A2(g127C),.A1(g6035C));
NAND2_X1 U_I7225C (.ZN(I7225C),.A2(I7223C),.A1(g1781C));
NAND2_X1 U_I11261C (.ZN(I11261C),.A2(g826C),.A1(g6775C));
NAND3_X1 U_g8843C (.ZN(g8843C),.A3(g8545C),.A2(g8757C),.A1(g8542C));
NAND2_X1 U_g2938C (.ZN(g2938C),.A2(I6111C),.A1(I6110C));
NAND2_X1 U_I4942C (.ZN(I4942C),.A2(I4941C),.A1(g396C));
NAND2_X1 U_g10394C (.ZN(g10394C),.A2(I15900C),.A1(I15899C));
NAND2_X1 U_g8549C (.ZN(g8549C),.A2(g8390C),.A1(g5527C));
NAND2_X1 U_g3070C (.ZN(g3070C),.A2(g1206C),.A1(g2016C));
NAND2_X1 U_I4954C (.ZN(I4954C),.A2(g327C),.A1(g401C));
NAND2_X1 U_I5023C (.ZN(I5023C),.A2(g1275C),.A1(g995C));
NAND2_X1 U_g10446C (.ZN(g10446C),.A2(g5350C),.A1(g10438C));
NAND2_X1 U_I16081C (.ZN(I16081C),.A2(I16079C),.A1(g10363C));
NAND2_X1 U_I8641C (.ZN(I8641C),.A2(I8640C),.A1(g4278C));
NAND2_X1 U_I6178C (.ZN(I6178C),.A2(I6176C),.A1(g197C));
NAND2_X1 U_I12075C (.ZN(I12075C),.A2(I12074C),.A1(g6015C));
NAND2_X1 U_I5127C (.ZN(I5127C),.A2(I5126C),.A1(g1386C));
NAND2_X1 U_I5451C (.ZN(I5451C),.A2(I5449C),.A1(g991C));
NAND2_X1 U_g4168C (.ZN(g4168C),.A2(I7323C),.A1(I7322C));
NAND2_X1 U_I6288C (.ZN(I6288C),.A2(I6287C),.A1(g2091C));
NAND2_X1 U_I8179C (.ZN(I8179C),.A2(I8178C),.A1(g3685C));
NAND2_X1 U_I4912C (.ZN(I4912C),.A2(I4910C),.A1(g318C));
NAND2_X1 U_I6805C (.ZN(I6805C),.A2(g471C),.A1(g3268C));
NAND3_X1 U_g3766C (.ZN(g3766C),.A3(g2493C),.A2(g3222C),.A1(g2439C));
NAND2_X1 U_g3087C (.ZN(g3087C),.A2(I6289C),.A1(I6288C));
NAND2_X1 U_I17486C (.ZN(I17486C),.A2(I17485C),.A1(g11233C));
NAND2_X1 U_I4929C (.ZN(I4929C),.A2(I4928C),.A1(g391C));
NAND2_X1 U_I15890C (.ZN(I15890C),.A2(g10285C),.A1(g853C));
NAND2_X1 U_I16331C (.ZN(I16331C),.A2(I16330C),.A1(g10387C));
NAND2_X1 U_I9575C (.ZN(I9575C),.A2(I9574C),.A1(g5608C));
NAND2_X1 U_I13887C (.ZN(I13887C),.A2(I13886C),.A1(g8267C));
NAND2_X1 U_g5308C (.ZN(g5308C),.A2(I8788C),.A1(I8787C));
NAND2_X1 U_I13529C (.ZN(I13529C),.A2(g8253C),.A1(g704C));
NAND2_X1 U_I6208C (.ZN(I6208C),.A2(I6207C),.A1(g5188C));
NAND2_X1 U_g5217C (.ZN(g5217C),.A2(I8642C),.A1(I8641C));
NAND2_X1 U_I5316C (.ZN(I5316C),.A2(I5315C),.A1(g1032C));
NAND2_X1 U_g2111C (.ZN(g2111C),.A2(I5007C),.A1(I5006C));
NAND2_X1 U_g10366C (.ZN(g10366C),.A2(g5392C),.A1(g10285C));
NAND2_X1 U_I5034C (.ZN(I5034C),.A2(g1019C),.A1(g1015C));
NAND2_X1 U_I13869C (.ZN(I13869C),.A2(I13867C),.A1(g1403C));
NAND2_X1 U_I13868C (.ZN(I13868C),.A2(I13867C),.A1(g8264C));
NAND2_X1 U_I15999C (.ZN(I15999C),.A2(FE_OFN247_g1771C),.A1(g10432C));
NAND2_X1 U_I13259C (.ZN(I13259C),.A2(I13258C),.A1(g1900C));
NAND4_X1 U_g3261C (.ZN(g3261C),.A4(g2202C),.A3(g2211C),.A2(g2222C),.A1(g2229C));
NAND2_X1 U_g10481C (.ZN(g10481C),.A2(I16074C),.A1(I16073C));
NAND2_X1 U_g2180C (.ZN(g2180C),.A2(I5137C),.A1(I5136C));
NAND3_X1 U_g4976C (.ZN(g4976C),.A3(g3807C),.A2(g4604C),.A1(g2310C));
NAND2_X1 U_g8506C (.ZN(g8506C),.A2(g8366C),.A1(g3475C));
NAND2_X1 U_g2380C (.ZN(g2380C),.A2(I5461C),.A1(I5460C));
NAND2_X1 U_I13258C (.ZN(I13258C),.A2(g8153C),.A1(g1900C));
NAND2_X1 U_I5013C (.ZN(I5013C),.A2(g1011C),.A1(g1007C));
NAND2_X1 U_g5196C (.ZN(g5196C),.A2(I8606C),.A1(I8605C));
NAND2_X1 U_I10930C (.ZN(I10930C),.A2(g5555C),.A1(g5863C));
NAND2_X1 U_I6770C (.ZN(I6770C),.A2(g382C),.A1(g3257C));
NAND2_X1 U_g11449C (.ZN(g11449C),.A2(I17402C),.A1(I17401C));
NAND2_X1 U_g11448C (.ZN(g11448C),.A2(I17395C),.A1(I17394C));
NAND2_X1 U_I15717C (.ZN(I15717C),.A2(I15716C),.A1(g10231C));
NAND2_X1 U_I5317C (.ZN(I5317C),.A2(I5315C),.A1(g1027C));
NAND2_X1 U_I14210C (.ZN(I14210C),.A2(I14209C),.A1(g8824C));
NAND2_X1 U_I17569C (.ZN(I17569C),.A2(I17567C),.A1(g1610C));
NAND2_X1 U_I13878C (.ZN(I13878C),.A2(I13876C),.A1(g1444C));
NAND2_X1 U_g8545C (.ZN(g8545C),.A2(g8390C),.A1(g3710C));
NAND2_X1 U_g2515C (.ZN(g2515C),.A2(I5606C),.A1(I5605C));
NAND2_X1 U_I14443C (.ZN(I14443C),.A2(I14442C),.A1(g8970C));
NAND2_X1 U_g7557C (.ZN(g7557C),.A2(I11997C),.A1(I11996C));
NAND2_X1 U_g8180C (.ZN(g8180C),.A2(I13091C),.A1(I13090C));
NAND2_X1 U_I14279C (.ZN(I14279C),.A2(I14277C),.A1(g1828C));
NAND2_X1 U_I17568C (.ZN(I17568C),.A2(I17567C),.A1(g11496C));
NAND2_X1 U_I13886C (.ZN(I13886C),.A2(g1440C),.A1(g8267C));
NAND2_X1 U_I7322C (.ZN(I7322C),.A2(I7321C),.A1(g3047C));
NAND2_X1 U_I6990C (.ZN(I6990C),.A2(I6988C),.A1(g986C));
NAND2_X1 U_I14278C (.ZN(I14278C),.A2(I14277C),.A1(g8847C));
NAND2_X1 U_I7033C (.ZN(I7033C),.A2(g1868C),.A1(g3089C));
NAND2_X1 U_I9006C (.ZN(I9006C),.A2(FE_OFN252_g1791C),.A1(g4492C));
NAND2_X1 U_g8507C (.ZN(g8507C),.A2(g8366C),.A1(g3738C));
NAND2_X1 U_I5460C (.ZN(I5460C),.A2(I5459C),.A1(g1240C));
NAND2_X1 U_g4588C (.ZN(g4588C),.A2(FE_OFN325_g18C),.A1(g3440C));
NAND2_X1 U_I4986C (.ZN(I4986C),.A2(I4985C),.A1(g999C));
NAND3_X1 U_g3247C (.ZN(g3247C),.A3(g2571C),.A2(g2564C),.A1(g1828C));
NAND2_X1 U_I8651C (.ZN(I8651C),.A2(I8650C),.A1(g4824C));
NAND2_X1 U_I13545C (.ZN(I13545C),.A2(I13544C),.A1(g713C));
NAND2_X1 U_g8628C (.ZN(g8628C),.A2(I13895C),.A1(I13894C));
NAND2_X1 U_I6138C (.ZN(I6138C),.A2(I6136C),.A1(g378C));
NAND2_X1 U_I12074C (.ZN(I12074C),.A2(g174C),.A1(g6015C));
NAND2_X1 U_g8630C (.ZN(g8630C),.A2(I13909C),.A1(I13908C));
NAND2_X1 U_I13078C (.ZN(I13078C),.A2(I13076C),.A1(g7963C));
NAND2_X1 U_I6109C (.ZN(I6109C),.A2(g1494C),.A1(g2205C));
NAND2_X1 U_g8300C (.ZN(g8300C),.A2(I13260C),.A1(I13259C));
NAND2_X1 U_I5501C (.ZN(I5501C),.A2(I5500C),.A1(g1255C));
NAND2_X1 U_I17586C (.ZN(I17586C),.A2(I17584C),.A1(g11515C));
NAND2_X1 U_I12092C (.ZN(I12092C),.A2(g1490C),.A1(g5810C));
NAND2_X1 U_I13901C (.ZN(I13901C),.A2(I13900C),.A1(g8261C));
NAND2_X1 U_I8795C (.ZN(I8795C),.A2(g1145C),.A1(g4672C));
NAND2_X1 U_I6201C (.ZN(I6201C),.A2(I6199C),.A1(g766C));
NAND2_X1 U_I14217C (.ZN(I14217C),.A2(I14216C),.A1(g8826C));
NAND2_X1 U_I9007C (.ZN(I9007C),.A2(I9006C),.A1(g4492C));
NAND2_X1 U_I13561C (.ZN(I13561C),.A2(I13559C),.A1(g8263C));
NAND2_X1 U_I15716C (.ZN(I15716C),.A2(g10229C),.A1(g10231C));
NAND2_X1 U_I6449C (.ZN(I6449C),.A2(I6447C),.A1(FE_OFN236_g1776C));
NAND2_X1 U_I13295C (.ZN(I13295C),.A2(I13293C),.A1(g8161C));
NAND2_X1 U_I4987C (.ZN(I4987C),.A2(I4985C),.A1(g1003C));
NAND2_X1 U_I6715C (.ZN(I6715C),.A2(I6714C),.A1(g2961C));
NAND2_X1 U_I17493C (.ZN(I17493C),.A2(I17492C),.A1(g11430C));
NAND2_X1 U_I12215C (.ZN(I12215C),.A2(I12214C),.A1(g7061C));
NAND2_X1 U_g2372C (.ZN(g2372C),.A2(I5451C),.A1(I5450C));
NAND2_X1 U_g7062C (.ZN(g7062C),.A2(I11263C),.A1(I11262C));
NAND2_X1 U_g2988C (.ZN(g2988C),.A2(I6226C),.A1(I6225C));
NAND2_X1 U_I13309C (.ZN(I13309C),.A2(I13307C),.A1(g617C));
NAND2_X1 U_g8839C (.ZN(g8839C),.A2(FE_OFN223_g4401C),.A1(g8603C));
NAND2_X1 U_g2555C (.ZN(g2555C),.A2(I5677C),.A1(I5676C));
NAND2_X1 U_g3662C (.ZN(g3662C),.A2(I6827C),.A1(I6826C));
NAND2_X1 U_I13308C (.ZN(I13308C),.A2(I13307C),.A1(g8190C));
NAND2_X1 U_g2792C (.ZN(g2792C),.A2(I5880C),.A1(I5879C));
NAND2_X1 U_g4117C (.ZN(g4117C),.A2(g3061C),.A1(g3041C));
NAND2_X1 U_I8543C (.ZN(I8543C),.A2(g486C),.A1(g4218C));
NAND2_X1 U_g11549C (.ZN(g11549C),.A2(I17586C),.A1(I17585C));
NAND2_X1 U_I6881C (.ZN(I6881C),.A2(I6879C),.A1(g1351C));
NAND2_X1 U_I12138C (.ZN(I12138C),.A2(I12136C),.A1(g131C));
NAND2_X1 U_I8729C (.ZN(I8729C),.A2(I8728C),.A1(g4605C));
NAND2_X1 U_I14216C (.ZN(I14216C),.A2(g605C),.A1(g8826C));
NAND2_X1 U_g10384C (.ZN(g10384C),.A2(I15872C),.A1(I15871C));
NAND2_X1 U_I13260C (.ZN(I13260C),.A2(I13258C),.A1(g8153C));
NAND2_X1 U_g2776C (.ZN(g2776C),.A2(I5867C),.A1(I5866C));
NAND2_X1 U_I8513C (.ZN(I8513C),.A2(g3513C),.A1(g4873C));
NAND2_X1 U_I13559C (.ZN(I13559C),.A2(g8263C),.A1(g722C));
NAND2_X1 U_I8178C (.ZN(I8178C),.A2(FE_OFN253_g1786C),.A1(g3685C));
NAND2_X1 U_g3631C (.ZN(g3631C),.A2(I6794C),.A1(I6793C));
NAND2_X1 U_I6487C (.ZN(I6487C),.A2(g1227C),.A1(g2306C));
NAND2_X1 U_I16080C (.ZN(I16080C),.A2(I16079C),.A1(g849C));
NAND2_X1 U_I13893C (.ZN(I13893C),.A2(g1436C),.A1(g8266C));
NAND2_X1 U_I12115C (.ZN(I12115C),.A2(I12113C),.A1(g162C));
NAND2_X1 U_I6748C (.ZN(I6748C),.A2(I6746C),.A1(g1453C));
NAND2_X1 U_I13544C (.ZN(I13544C),.A2(g8259C),.A1(g713C));
NAND2_X1 U_I5484C (.ZN(I5484C),.A2(g1011C),.A1(g1250C));
NAND2_X1 U_I4928C (.ZN(I4928C),.A2(g321C),.A1(g391C));
NAND2_X1 U_I6226C (.ZN(I6226C),.A2(I6224C),.A1(g1346C));
NAND2_X1 U_I8805C (.ZN(I8805C),.A2(I8803C),.A1(g1113C));
NAND2_X1 U_I4930C (.ZN(I4930C),.A2(I4928C),.A1(g321C));
NAND2_X1 U_I15880C (.ZN(I15880C),.A2(I15878C),.A1(FE_OFN251_g1801C));
NAND2_X1 U_I14265C (.ZN(I14265C),.A2(I14263C),.A1(g1814C));
NAND2_X1 U_I16031C (.ZN(I16031C),.A2(I16030C),.A1(g829C));
NAND2_X1 U_g3585C (.ZN(g3585C),.A2(I6748C),.A1(I6747C));
NAND4_X1 U_g3041C (.ZN(g3041C),.A4(g2382C),.A3(g2374C),.A2(g2399C),.A1(g2364C));
NAND2_X1 U_g8933C (.ZN(g8933C),.A2(I14272C),.A1(I14271C));
NAND2_X1 U_I16330C (.ZN(I16330C),.A2(g4997C),.A1(g10387C));
NAND2_X1 U_I13267C (.ZN(I13267C),.A2(I13265C),.A1(g8154C));
NAND2_X1 U_I13294C (.ZN(I13294C),.A2(I13293C),.A1(g1882C));
NAND2_X1 U_g10231C (.ZN(g10231C),.A2(I15617C),.A1(I15616C));
NAND2_X1 U_I14442C (.ZN(I14442C),.A2(g1834C),.A1(g8970C));
NAND2_X1 U_I6793C (.ZN(I6793C),.A2(I6792C),.A1(g2959C));
NAND2_X1 U_I4966C (.ZN(I4966C),.A2(I4964C),.A1(g330C));
NAND2_X1 U_I8752C (.ZN(I8752C),.A2(I8750C),.A1(g1125C));
NAND2_X1 U_I15432C (.ZN(I15432C),.A2(I15430C),.A1(g9995C));
NAND2_X1 U_I12214C (.ZN(I12214C),.A2(g2518C),.A1(g7061C));
NAND2_X1 U_g10511C (.ZN(g10511C),.A2(g6032C),.A1(g10438C));
NAND2_X1 U_g3011C (.ZN(g3011C),.A2(g2382C),.A1(g591C));
NAND2_X1 U_g5103C (.ZN(g5103C),.A2(I8481C),.A1(I8480C));
NAND2_X1 U_I16087C (.ZN(I16087C),.A2(I16086C),.A1(g861C));
NAND2_X1 U_g3734C (.ZN(g3734C),.A2(g599C),.A1(g3039C));
NAND2_X1 U_I6664C (.ZN(I6664C),.A2(g2776C),.A1(g2792C));
NAND2_X1 U_g8882C (.ZN(g8882C),.A2(I14218C),.A1(I14217C));
NAND2_X1 U_I4955C (.ZN(I4955C),.A2(I4954C),.A1(g401C));
NAND2_X1 U_I8786C (.ZN(I8786C),.A2(g1141C),.A1(g4639C));
NAND3_X1 U_g3992C (.ZN(g3992C),.A3(g2990C),.A2(g2550C),.A1(g2571C));
NAND2_X1 U_g10480C (.ZN(g10480C),.A2(I16067C),.A1(I16066C));
NAND2_X1 U_I11915C (.ZN(I11915C),.A2(I11914C),.A1(g5803C));
NAND2_X1 U_I8770C (.ZN(I8770C),.A2(g1133C),.A1(g4619C));
NAND2_X1 U_I5516C (.ZN(I5516C),.A2(g1019C),.A1(g1260C));
NAND2_X1 U_g8541C (.ZN(g8541C),.A2(g8390C),.A1(g4001C));
NAND2_X1 U_I6188C (.ZN(I6188C),.A2(I6186C),.A1(g466C));
NAND2_X1 U_g5147C (.ZN(g5147C),.A2(I8545C),.A1(I8544C));
NAND3_X1 U_g8744C (.ZN(g8744C),.A3(I9273C),.A2(g46C),.A1(g8617C));
NAND2_X1 U_I5892C (.ZN(I5892C),.A2(I5891C),.A1(g750C));
NAND2_X1 U_g8558C (.ZN(g8558C),.A2(I13767C),.A1(I13766C));
NAND2_X1 U_I15258C (.ZN(I15258C),.A2(I15256C),.A1(g9968C));
NAND2_X1 U_I13266C (.ZN(I13266C),.A2(I13265C),.A1(g1909C));
NAND2_X1 U_I8787C (.ZN(I8787C),.A2(I8786C),.A1(g4639C));
NAND2_X1 U_I6826C (.ZN(I6826C),.A2(I6825C),.A1(g3281C));
NAND2_X1 U_I17283C (.ZN(I17283C),.A2(I17281C),.A1(g11219C));
NAND3_X1 U_g5013C (.ZN(g5013C),.A3(g3205C),.A2(g3247C),.A1(g4749C));
NAND2_X1 U_I17492C (.ZN(I17492C),.A2(g3623C),.A1(g11430C));
NAND2_X1 U_g8511C (.ZN(g8511C),.A2(g8366C),.A1(g5277C));
NAND2_X1 U_I16079C (.ZN(I16079C),.A2(g10363C),.A1(g849C));
NAND2_X1 U_I5035C (.ZN(I5035C),.A2(I5034C),.A1(g1015C));
NAND2_X1 U_I5517C (.ZN(I5517C),.A2(I5516C),.A1(g1260C));
NAND2_X1 U_I7223C (.ZN(I7223C),.A2(g1781C),.A1(g2981C));
NAND2_X1 U_I16086C (.ZN(I16086C),.A2(g10430C),.A1(g861C));
NAND2_X1 U_g5317C (.ZN(g5317C),.A2(I8797C),.A1(I8796C));
NAND2_X1 U_I15879C (.ZN(I15879C),.A2(I15878C),.A1(g10359C));
NAND2_X1 U_I15878C (.ZN(I15878C),.A2(FE_OFN251_g1801C),.A1(g10359C));
NAND2_X1 U_I12114C (.ZN(I12114C),.A2(I12113C),.A1(g6002C));
NAND2_X1 U_I12107C (.ZN(I12107C),.A2(I12106C),.A1(g6042C));
NAND2_X1 U_g2500C (.ZN(g2500C),.A2(g182C),.A1(g178C));
NAND2_X1 U_I15994C (.ZN(I15994C),.A2(I15992C),.A1(g2677C));
NAND4_X1 U_g7934C (.ZN(g7934C),.A4(g7550C),.A3(FE_OFN91_g2172C),.A2(FE_OFN80_g2175C),.A1(g6941C));
NAND2_X1 U_g10469C (.ZN(g10469C),.A2(g5999C),.A1(g10430C));
NAND2_X1 U_I14264C (.ZN(I14264C),.A2(I14263C),.A1(g8843C));
NAND2_X1 U_I6448C (.ZN(I6448C),.A2(I6447C),.A1(g2264C));
NAND2_X1 U_I13285C (.ZN(I13285C),.A2(I13283C),.A1(g8159C));
NAND2_X1 U_g10468C (.ZN(g10468C),.A2(I16001C),.A1(I16000C));
NAND2_X1 U_I6827C (.ZN(I6827C),.A2(I6825C),.A1(g770C));
NAND2_X1 U_g8623C (.ZN(g8623C),.A2(I13878C),.A1(I13877C));
NAND2_X1 U_I13900C (.ZN(I13900C),.A2(g1428C),.A1(g8261C));
NAND2_X1 U_g2795C (.ZN(g2795C),.A2(I5893C),.A1(I5892C));
NAND2_X1 U_I8575C (.ZN(I8575C),.A2(g496C),.A1(g4234C));
NAND2_X1 U_I14209C (.ZN(I14209C),.A2(g599C),.A1(g8824C));
NAND2_X1 U_I13560C (.ZN(I13560C),.A2(I13559C),.A1(g722C));
NAND2_X1 U_I8715C (.ZN(I8715C),.A2(g4052C),.A1(g4601C));
NAND2_X1 U_I8604C (.ZN(I8604C),.A2(g506C),.A1(g4259C));
NAND2_X1 U_I16017C (.ZN(I16017C),.A2(I16015C),.A1(g1781C));
NAND2_X1 U_I4941C (.ZN(I4941C),.A2(g324C),.A1(g396C));
NAND2_X1 U_g2205C (.ZN(g2205C),.A2(I5166C),.A1(I5165C));
NAND3_X1 U_g3753C (.ZN(g3753C),.A3(g2800C),.A2(g2364C),.A1(g2382C));
NAND2_X1 U_I6467C (.ZN(I6467C),.A2(g2479C),.A1(g23C));
NAND2_X1 U_I14614C (.ZN(I14614C),.A2(I14612C),.A1(g611C));
NAND2_X1 U_g2104C (.ZN(g2104C),.A2(I4966C),.A1(I4965C));
NAND2_X1 U_g2099C (.ZN(g2099C),.A2(I4943C),.A1(I4942C));
NAND2_X1 U_I16023C (.ZN(I16023C),.A2(FE_OFN253_g1786C),.A1(g10438C));
NAND2_X1 U_g10479C (.ZN(g10479C),.A2(I16060C),.A1(I16059C));
NAND3_X1 U_g8737C (.ZN(g8737C),.A3(g8688C),.A2(FE_OFN200_g4921C),.A1(g1975C));
NAND2_X1 U_g5942C (.ZN(g5942C),.A2(I9576C),.A1(I9575C));
NAND2_X1 U_g10478C (.ZN(g10478C),.A2(I16053C),.A1(I16052C));
NAND2_X1 U_I12004C (.ZN(I12004C),.A2(I12002C),.A1(g153C));
NAND2_X1 U_I4911C (.ZN(I4911C),.A2(I4910C),.A1(g386C));
NAND2_X1 U_I11914C (.ZN(I11914C),.A2(g1494C),.A1(g5803C));
NAND2_X1 U_g7960C (.ZN(g7960C),.A2(g5573C),.A1(g7409C));
NAND2_X1 U_I5295C (.ZN(I5295C),.A2(g798C),.A1(g794C));
NAND2_X1 U_I12106C (.ZN(I12106C),.A2(g135C),.A1(g6042C));
NAND2_X1 U_I8728C (.ZN(I8728C),.A2(g1117C),.A1(g4605C));
NAND2_X1 U_g3681C (.ZN(g3681C),.A2(I6838C),.A1(I6837C));
NAND2_X1 U_I11907C (.ZN(I11907C),.A2(g1474C),.A1(g5838C));
NAND2_X1 U_I13907C (.ZN(I13907C),.A2(g1432C),.A1(g8265C));
NAND2_X1 U_I8730C (.ZN(I8730C),.A2(I8728C),.A1(g1117C));
NAND2_X1 U_g8551C (.ZN(g8551C),.A2(g8390C),.A1(g3967C));
NAND2_X1 U_I4980C (.ZN(I4980C),.A2(I4978C),.A1(g333C));
NAND2_X1 U_g2961C (.ZN(g2961C),.A2(I6178C),.A1(I6177C));
NAND2_X1 U_g6019C (.ZN(g6019C),.A2(FE_OFN200_g4921C),.A1(g617C));
NAND2_X1 U_I16016C (.ZN(I16016C),.A2(I16015C),.A1(g10441C));
NAND2_X1 U_I11935C (.ZN(I11935C),.A2(g1458C),.A1(g5857C));
NAND2_X1 U_I8678C (.ZN(I8678C),.A2(I8676C),.A1(g1027C));
NAND2_X1 U_I17051C (.ZN(I17051C),.A2(g11249C),.A1(g10923C));
NAND2_X1 U_g4482C (.ZN(g4482C),.A2(I7865C),.A1(I7864C));
NAND2_X1 U_g7592C (.ZN(g7592C),.A2(I12108C),.A1(I12107C));
NAND2_X1 U_g3460C (.ZN(g3460C),.A2(I6666C),.A1(I6665C));
NAND4_X1 U_g7932C (.ZN(g7932C),.A4(FE_OFN96_g2169C),.A3(FE_OFN91_g2172C),.A2(FE_OFN80_g2175C),.A1(g6941C));
NAND2_X1 U_g7624C (.ZN(g7624C),.A2(I12216C),.A1(I12215C));
NAND4_X1 U_g7953C (.ZN(g7953C),.A4(g7550C),.A3(g7562C),.A2(g7574C),.A1(g6941C));
NAND2_X1 U_g8414C (.ZN(g8414C),.A2(I13554C),.A1(I13553C));
NAND2_X1 U_I6168C (.ZN(I6168C),.A2(I6166C),.A1(g153C));
NAND2_X1 U_I5229C (.ZN(I5229C),.A2(g148C),.A1(g182C));
NAND2_X1 U_I6772C (.ZN(I6772C),.A2(I6770C),.A1(g382C));
NAND2_X1 U_I16030C (.ZN(I16030C),.A2(g10430C),.A1(g829C));
NAND2_X1 U_I13284C (.ZN(I13284C),.A2(I13283C),.A1(g1927C));
NAND2_X1 U_I16065C (.ZN(I16065C),.A2(FE_OFN237_g1806C),.A1(g10428C));
NAND2_X1 U_g2947C (.ZN(g2947C),.A2(I6138C),.A1(I6137C));
NAND2_X1 U_I7321C (.ZN(I7321C),.A2(g1231C),.A1(g3047C));
NAND2_X1 U_g2437C (.ZN(g2437C),.A2(I5530C),.A1(I5529C));
NAND2_X1 U_g2102C (.ZN(g2102C),.A2(I4956C),.A1(I4955C));
NAND2_X1 U_I17282C (.ZN(I17282C),.A2(I17281C),.A1(g11221C));
NAND2_X1 U_I5620C (.ZN(I5620C),.A2(I5618C),.A1(FE_OFN247_g1771C));
NAND2_X1 U_I8664C (.ZN(I8664C),.A2(I8662C),.A1(g476C));
NAND2_X1 U_g7524C (.ZN(g7524C),.A2(I11916C),.A1(I11915C));
NAND2_X1 U_g7717C (.ZN(g7717C),.A2(g1950C),.A1(g6863C));
NAND2_X1 U_I16467C (.ZN(I16467C),.A2(g10518C),.A1(g10716C));
NAND2_X1 U_I4972C (.ZN(I4972C),.A2(I4971C),.A1(g991C));
NAND2_X1 U_I13554C (.ZN(I13554C),.A2(I13552C),.A1(g8262C));
NAND2_X1 U_I16037C (.ZN(I16037C),.A2(FE_OFN252_g1791C),.A1(g10363C));
NAND2_X1 U_g8302C (.ZN(g8302C),.A2(I13274C),.A1(I13273C));
NAND2_X1 U_I4943C (.ZN(I4943C),.A2(I4941C),.A1(g324C));
NAND2_X1 U_I5485C (.ZN(I5485C),.A2(I5484C),.A1(g1250C));
NAND2_X1 U_g5527C (.ZN(g5527C),.A2(g4749C),.A1(g3978C));
NAND2_X1 U_I10509C (.ZN(I10509C),.A2(I10507C),.A1(g786C));
NAND2_X1 U_g7599C (.ZN(g7599C),.A2(I12145C),.A1(I12144C));
NAND2_X1 U_I10508C (.ZN(I10508C),.A2(I10507C),.A1(g6221C));
NAND2_X1 U_I6126C (.ZN(I6126C),.A2(I6124C),.A1(g1419C));
NAND2_X1 U_I8671C (.ZN(I8671C),.A2(I8669C),.A1(g814C));
NAND2_X1 U_I6760C (.ZN(I6760C),.A2(g1448C),.A1(g2943C));
NAND2_X1 U_g3626C (.ZN(g3626C),.A2(I6779C),.A1(I6778C));
NAND2_X1 U_I11973C (.ZN(I11973C),.A2(g1462C),.A1(g5852C));
NAND2_X1 U_g2389C (.ZN(g2389C),.A2(I5470C),.A1(I5469C));
NAND2_X1 U_I15617C (.ZN(I15617C),.A2(I15615C),.A1(g10153C));
NAND2_X1 U_g5277C (.ZN(g5277C),.A2(g4538C),.A1(g3734C));
NAND2_X1 U_I5005C (.ZN(I5005C),.A2(g312C),.A1(g421C));
NAND2_X1 U_I6779C (.ZN(I6779C),.A2(I6777C),.A1(g650C));
NAND2_X1 U_I6665C (.ZN(I6665C),.A2(I6664C),.A1(g2792C));
NAND2_X1 U_I8589C (.ZN(I8589C),.A2(g501C),.A1(g4251C));
NAND2_X1 U_g8412C (.ZN(g8412C),.A2(I13546C),.A1(I13545C));
NAND2_X1 U_g2963C (.ZN(g2963C),.A2(I6188C),.A1(I6187C));
NAND2_X1 U_I12045C (.ZN(I12045C),.A2(g1486C),.A1(g5814C));
NAND2_X1 U_I16053C (.ZN(I16053C),.A2(I16051C),.A1(g10434C));
NAND2_X1 U_g2109C (.ZN(g2109C),.A2(I4997C),.A1(I4996C));
NAND2_X1 U_g11418C (.ZN(g11418C),.A2(I17307C),.A1(I17306C));
NAND2_X1 U_I13539C (.ZN(I13539C),.A2(I13537C),.A1(g8157C));
NAND2_X1 U_g10475C (.ZN(g10475C),.A2(I16032C),.A1(I16031C));
NAND2_X1 U_I5324C (.ZN(I5324C),.A2(I5323C),.A1(g1336C));
NAND2_X1 U_I13538C (.ZN(I13538C),.A2(I13537C),.A1(g658C));
NAND2_X1 U_I5469C (.ZN(I5469C),.A2(I5468C),.A1(g1245C));
NAND2_X1 U_I5540C (.ZN(I5540C),.A2(I5538C),.A1(g1023C));
NAND2_X1 U_I17505C (.ZN(I17505C),.A2(I17503C),.A1(g5269C));
NAND2_X1 U_I11241C (.ZN(I11241C),.A2(g790C),.A1(g6760C));
NAND2_X1 U_I8803C (.ZN(I8803C),.A2(g1113C),.A1(g4677C));
NAND2_X1 U_I12061C (.ZN(I12061C),.A2(I12060C),.A1(g5824C));
NAND2_X1 U_I8780C (.ZN(I8780C),.A2(I8778C),.A1(g1137C));
NAND3_X1 U_g8745C (.ZN(g8745C),.A3(I9265C),.A2(g47C),.A1(g8617C));
NAND2_X1 U_I4979C (.ZN(I4979C),.A2(I4978C),.A1(g411C));
NAND2_X1 U_g8109C (.ZN(g8109C),.A2(I11360C),.A1(g48C));
NAND2_X1 U_g8309C (.ZN(g8309C),.A2(I13309C),.A1(I13308C));
NAND2_X1 U_g6758C (.ZN(g6758C),.A2(I10771C),.A1(I10770C));
NAND2_X1 U_I16009C (.ZN(I16009C),.A2(I16007C),.A1(FE_OFN236_g1776C));
NAND2_X1 U_I15616C (.ZN(I15616C),.A2(I15615C),.A1(g10043C));
NAND2_X1 U_I8662C (.ZN(I8662C),.A2(g476C),.A1(g4286C));
NAND2_X1 U_I16008C (.ZN(I16008C),.A2(I16007C),.A1(g10434C));
NAND2_X1 U_I13515C (.ZN(I13515C),.A2(I13513C),.A1(g8248C));
NAND2_X1 U_I13991C (.ZN(I13991C),.A2(I13990C),.A1(g622C));
NAND2_X1 U_g11276C (.ZN(g11276C),.A2(I17053C),.A1(I17052C));
NAND2_X1 U_I15900C (.ZN(I15900C),.A2(I15898C),.A1(g10359C));
NAND2_X1 U_g2419C (.ZN(g2419C),.A2(I5502C),.A1(I5501C));
NAND2_X1 U_I16074C (.ZN(I16074C),.A2(I16072C),.A1(g10438C));
NAND2_X1 U_I10769C (.ZN(I10769C),.A2(FE_OFN251_g1801C),.A1(g5944C));
NAND2_X1 U_I7323C (.ZN(I7323C),.A2(I7321C),.A1(g1231C));
NAND2_X1 U_g7978C (.ZN(g7978C),.A2(g736C),.A1(g7697C));
NAND2_X1 U_I7875C (.ZN(I7875C),.A2(g810C),.A1(g4109C));
NAND2_X1 U_I8562C (.ZN(I8562C),.A2(I8561C),.A1(g4227C));
NAND2_X1 U_I15892C (.ZN(I15892C),.A2(I15890C),.A1(g10285C));
NAND2_X1 U_g3771C (.ZN(g3771C),.A2(I6990C),.A1(I6989C));
NAND2_X1 U_I8605C (.ZN(I8605C),.A2(I8604C),.A1(g4259C));
NAND2_X1 U_g10153C (.ZN(g10153C),.A2(I15453C),.A1(I15452C));
NAND2_X1 U_g5295C (.ZN(g5295C),.A2(I8763C),.A1(I8762C));
NAND2_X1 U_I8751C (.ZN(I8751C),.A2(I8750C),.A1(g4613C));
NAND2_X1 U_I15907C (.ZN(I15907C),.A2(I15906C),.A1(g6899C));
NAND2_X1 U_I5136C (.ZN(I5136C),.A2(I5135C),.A1(g521C));
NAND2_X1 U_I11263C (.ZN(I11263C),.A2(I11261C),.A1(g826C));
NAND2_X1 U_I14204C (.ZN(I14204C),.A2(I14202C),.A1(g591C));
NAND2_X1 U_g8881C (.ZN(g8881C),.A2(I14211C),.A1(I14210C));
NAND2_X1 U_g2105C (.ZN(g2105C),.A2(I4973C),.A1(I4972C));
NAND3_X1 U_g5557C (.ZN(g5557C),.A3(g3011C),.A2(g3071C),.A1(g4538C));
NAND2_X1 U_I5230C (.ZN(I5230C),.A2(I5229C),.A1(g182C));
NAND2_X1 U_I8669C (.ZN(I8669C),.A2(g814C),.A1(g4831C));
NAND2_X1 U_g10474C (.ZN(g10474C),.A2(I16025C),.A1(I16024C));
NAND2_X1 U_I8772C (.ZN(I8772C),.A2(I8770C),.A1(g1133C));
NAND2_X1 U_g2445C (.ZN(g2445C),.A2(I5540C),.A1(I5539C));
NAND2_X1 U_g8006C (.ZN(g8006C),.A2(g7717C),.A1(g5552C));
NAND2_X1 U_I10932C (.ZN(I10932C),.A2(I10930C),.A1(g5555C));
NAND2_X1 U_I17504C (.ZN(I17504C),.A2(I17503C),.A1(g11430C));
NAND2_X1 U_I5137C (.ZN(I5137C),.A2(I5135C),.A1(g525C));
NAND2_X1 U_g8305C (.ZN(g8305C),.A2(I13285C),.A1(I13284C));
NAND2_X1 U_I5891C (.ZN(I5891C),.A2(g2057C),.A1(g750C));
NAND2_X1 U_I13273C (.ZN(I13273C),.A2(I13272C),.A1(g1918C));
NAND2_X1 U_I8480C (.ZN(I8480C),.A2(I8479C),.A1(g4455C));
NAND2_X2 U_g4144C (.ZN(g4144C),.A2(g109C),.A1(g2160C));
NAND2_X1 U_I15906C (.ZN(I15906C),.A2(g10302C),.A1(g6899C));
NAND2_X1 U_I5342C (.ZN(I5342C),.A2(I5341C),.A1(g315C));
NAND2_X1 U_I13514C (.ZN(I13514C),.A2(I13513C),.A1(g686C));
NAND2_X1 U_g8407C (.ZN(g8407C),.A2(I13523C),.A1(I13522C));
NAND2_X1 U_g4088C (.ZN(g4088C),.A2(I7225C),.A1(I7224C));
NAND2_X1 U_g4488C (.ZN(g4488C),.A2(I7877C),.A1(I7876C));
NAND2_X1 U_g7598C (.ZN(g7598C),.A2(I12138C),.A1(I12137C));
NAND3_X1 U_g3222C (.ZN(g3222C),.A3(g1834C),.A2(g1814C),.A1(g2557C));
NAND2_X1 U_I16052C (.ZN(I16052C),.A2(I16051C),.A1(g837C));
NAND2_X1 U_I12127C (.ZN(I12127C),.A2(I12126C),.A1(g6026C));
NAND2_X1 U_g10483C (.ZN(g10483C),.A2(I16088C),.A1(I16087C));
NAND2_X1 U_g8415C (.ZN(g8415C),.A2(I13561C),.A1(I13560C));
NAND2_X1 U_g11415C (.ZN(g11415C),.A2(I17290C),.A1(I17289C));
NAND2_X1 U_g6573C (.ZN(g6573C),.A2(I10509C),.A1(I10508C));
NAND2_X1 U_I5676C (.ZN(I5676C),.A2(I5675C),.A1(g1218C));
NAND2_X1 U_I6778C (.ZN(I6778C),.A2(I6777C),.A1(g2892C));
NAND2_X1 U_g9413C (.ZN(g9413C),.A2(I14614C),.A1(I14613C));
NAND2_X1 U_I8779C (.ZN(I8779C),.A2(I8778C),.A1(g4630C));
NAND2_X1 U_I5592C (.ZN(I5592C),.A2(I5591C),.A1(g1696C));
NAND4_X1 U_g8502C (.ZN(g8502C),.A4(g8366C),.A3(g591C),.A2(g605C),.A1(g2382C));
NAND2_X1 U_I15609C (.ZN(I15609C),.A2(I15607C),.A1(g10144C));
NAND2_X1 U_I15608C (.ZN(I15608C),.A2(I15607C),.A1(g10149C));
NAND3_X1 U_g3071C (.ZN(g3071C),.A3(g2382C),.A2(g2374C),.A1(g605C));
NAND2_X1 U_g10509C (.ZN(g10509C),.A2(g6023C),.A1(g10436C));
NAND2_X1 U_I17461C (.ZN(I17461C),.A2(I17459C),.A1(g11448C));
NAND2_X1 U_I13506C (.ZN(I13506C),.A2(I13504C),.A1(g8247C));
NAND2_X1 U_I5468C (.ZN(I5468C),.A2(g999C),.A1(g1245C));
NAND2_X1 U_g5219C (.ZN(g5219C),.A2(I8652C),.A1(I8651C));
NAND2_X1 U_I5677C (.ZN(I5677C),.A2(I5675C),.A1(g1223C));
NAND3_X1 U_g8826C (.ZN(g8826C),.A3(g8648C),.A2(g8737C),.A1(g8512C));
NAND2_X1 U_I17393C (.ZN(I17393C),.A2(g11414C),.A1(g11415C));
NAND2_X1 U_I5866C (.ZN(I5866C),.A2(I5865C),.A1(g2107C));
NAND2_X1 U_I12126C (.ZN(I12126C),.A2(g170C),.A1(g6026C));
NAND2_X1 U_I4978C (.ZN(I4978C),.A2(g333C),.A1(g411C));
NAND2_X1 U_g7587C (.ZN(g7587C),.A2(I12087C),.A1(I12086C));
NAND2_X1 U_g5286C (.ZN(g5286C),.A2(I8752C),.A1(I8751C));
NAND2_X1 U_g8308C (.ZN(g8308C),.A2(I13302C),.A1(I13301C));
NAND2_X1 U_I7864C (.ZN(I7864C),.A2(I7863C),.A1(g4099C));
NAND2_X1 U_I11981C (.ZN(I11981C),.A2(I11980C),.A1(g5820C));
NAND2_X1 U_I12060C (.ZN(I12060C),.A2(g1478C),.A1(g5824C));
NAND2_X1 U_g5225C (.ZN(g5225C),.A2(I8664C),.A1(I8663C));
NAND2_X1 U_g11538C (.ZN(g11538C),.A2(I17569C),.A1(I17568C));
NAND2_X1 U_I13767C (.ZN(I13767C),.A2(I13765C),.A1(g8417C));
NAND2_X1 U_g10396C (.ZN(g10396C),.A2(I15908C),.A1(I15907C));
NAND2_X1 U_I11262C (.ZN(I11262C),.A2(I11261C),.A1(g6775C));
NAND2_X1 U_I13990C (.ZN(I13990C),.A2(g8688C),.A1(g622C));
NAND2_X1 U_I6224C (.ZN(I6224C),.A2(g1346C),.A1(g2544C));
NAND2_X1 U_I5867C (.ZN(I5867C),.A2(I5865C),.A1(g2105C));
NAND2_X1 U_g2493C (.ZN(g2493C),.A2(g1840C),.A1(g1834C));
NAND2_X1 U_I5893C (.ZN(I5893C),.A2(I5891C),.A1(g2057C));
NAND3_X1 U_g3062C (.ZN(g3062C),.A3(g611C),.A2(g591C),.A1(g2369C));
NAND2_X1 U_I13521C (.ZN(I13521C),.A2(g8249C),.A1(g695C));
NAND2_X1 U_I5186C (.ZN(I5186C),.A2(I5184C),.A1(g1515C));
NAND2_X1 U_I6771C (.ZN(I6771C),.A2(I6770C),.A1(g3257C));
NAND2_X1 U_I5325C (.ZN(I5325C),.A2(I5323C),.A1(g1341C));
NAND2_X1 U_I17459C (.ZN(I17459C),.A2(g11448C),.A1(g11449C));
NAND2_X1 U_I9557C (.ZN(I9557C),.A2(g782C),.A1(g5598C));
NAND2_X1 U_g11414C (.ZN(g11414C),.A2(I17283C),.A1(I17282C));
NAND2_X1 U_I12067C (.ZN(I12067C),.A2(g139C),.A1(g6045C));
NAND2_X1 U_I12094C (.ZN(I12094C),.A2(I12092C),.A1(g1490C));
NAND2_X1 U_I4964C (.ZN(I4964C),.A2(g330C),.A1(g406C));
NAND2_X1 U_I13272C (.ZN(I13272C),.A2(g8158C),.A1(g1918C));
NAND2_X1 U_I9948C (.ZN(I9948C),.A2(I9946C),.A1(g1796C));
NAND2_X1 U_g10302C (.ZN(g10302C),.A2(I15718C),.A1(I15717C));
NAND2_X1 U_I16332C (.ZN(I16332C),.A2(I16330C),.A1(g4997C));
NAND2_X1 U_I5106C (.ZN(I5106C),.A2(I5104C),.A1(g435C));
NAND2_X1 U_g8847C (.ZN(g8847C),.A2(g8683C),.A1(g8551C));
NAND2_X1 U_g2257C (.ZN(g2257C),.A2(I5284C),.A1(I5283C));
NAND2_X1 U_I12019C (.ZN(I12019C),.A2(g166C),.A1(g6049C));
NAND2_X1 U_I15441C (.ZN(I15441C),.A2(g10007C),.A1(g10013C));
NAND2_X1 U_I11997C (.ZN(I11997C),.A2(I11995C),.A1(g127C));
NAND2_X1 U_I8739C (.ZN(I8739C),.A2(I8738C),.A1(g4607C));
NAND2_X1 U_I5461C (.ZN(I5461C),.A2(I5459C),.A1(g1003C));
NAND2_X1 U_I13766C (.ZN(I13766C),.A2(I13765C),.A1(g731C));
NAND2_X1 U_I8479C (.ZN(I8479C),.A2(g3530C),.A1(g4455C));
NAND2_X1 U_I17295C (.ZN(I17295C),.A2(g11227C),.A1(g11229C));
NAND2_X1 U_I14271C (.ZN(I14271C),.A2(I14270C),.A1(g8840C));
NAND2_X1 U_I4971C (.ZN(I4971C),.A2(g995C),.A1(g991C));
NAND2_X1 U_g8301C (.ZN(g8301C),.A2(I13267C),.A1(I13266C));
NAND2_X1 U_I6110C (.ZN(I6110C),.A2(I6109C),.A1(g2205C));
NAND2_X1 U_g10482C (.ZN(g10482C),.A2(I16081C),.A1(I16080C));
NAND2_X1 U_g10779C (.ZN(g10779C),.A2(I16469C),.A1(I16468C));
NAND2_X1 U_I6762C (.ZN(I6762C),.A2(I6760C),.A1(g1448C));
NAND2_X1 U_I17289C (.ZN(I17289C),.A2(I17288C),.A1(g11225C));
NAND2_X1 U_I5315C (.ZN(I5315C),.A2(g1027C),.A1(g1032C));
NAND2_X1 U_I17288C (.ZN(I17288C),.A2(g11223C),.A1(g11225C));
NAND2_X1 U_I13859C (.ZN(I13859C),.A2(I13857C),.A1(g1448C));
NAND2_X1 U_g7548C (.ZN(g7548C),.A2(I11982C),.A1(I11981C));
NAND2_X1 U_I13858C (.ZN(I13858C),.A2(I13857C),.A1(g8270C));
NAND2_X1 U_I11996C (.ZN(I11996C),.A2(I11995C),.A1(g6035C));
NAND3_X1 U_g8743C (.ZN(g8743C),.A3(I9265C),.A2(I9273C),.A1(g8617C));
NAND2_X1 U_I5880C (.ZN(I5880C),.A2(I5878C),.A1(g2115C));
NAND2_X1 U_g10513C (.ZN(g10513C),.A2(g5345C),.A1(g10441C));
NAND2_X1 U_g8411C (.ZN(g8411C),.A2(I13539C),.A1(I13538C));
NAND2_X1 U_I8626C (.ZN(I8626C),.A2(I8624C),.A1(g511C));
NAND2_X1 U_g10505C (.ZN(g10505C),.A2(g5938C),.A1(g10432C));
NAND2_X1 U_I5612C (.ZN(I5612C),.A2(I5611C),.A1(g1280C));
NAND2_X1 U_g4821C (.ZN(g4821C),.A2(I8180C),.A1(I8179C));
NAND2_X1 U_I12076C (.ZN(I12076C),.A2(I12074C),.A1(g174C));
NAND2_X1 U_I12085C (.ZN(I12085C),.A2(g1470C),.A1(g5842C));
NAND2_X1 U_g7567C (.ZN(g7567C),.A2(I12021C),.A1(I12020C));
NAND2_X1 U_I5128C (.ZN(I5128C),.A2(I5126C),.A1(g1389C));
NAND2_X1 U_I6489C (.ZN(I6489C),.A2(I6487C),.A1(g1227C));
NAND2_X1 U_g7593C (.ZN(g7593C),.A2(I12115C),.A1(I12114C));
NAND2_X1 U_I8778C (.ZN(I8778C),.A2(g1137C),.A1(g4630C));
NAND2_X1 U_g10149C (.ZN(g10149C),.A2(I15443C),.A1(I15442C));
NAND2_X1 U_I13902C (.ZN(I13902C),.A2(I13900C),.A1(g1428C));
NAND2_X1 U_I13301C (.ZN(I13301C),.A2(I13300C),.A1(g1936C));
NAND2_X1 U_g3215C (.ZN(g3215C),.A2(g1822C),.A1(g2564C));
NAND4_X1 U_g7996C (.ZN(g7996C),.A4(FE_OFN96_g2169C),.A3(g7562C),.A2(g7574C),.A1(FE_OFN88_g2178C));
NAND2_X1 U_I4985C (.ZN(I4985C),.A2(g1003C),.A1(g999C));
NAND2_X1 U_I14444C (.ZN(I14444C),.A2(I14442C),.A1(g1834C));
NAND4_X1 U_g8000C (.ZN(g8000C),.A4(g7550C),.A3(g7562C),.A2(g7574C),.A1(FE_OFN88_g2178C));
NAND2_X1 U_I5166C (.ZN(I5166C),.A2(I5164C),.A1(g1499C));
NAND2_X1 U_I17460C (.ZN(I17460C),.A2(I17459C),.A1(g11449C));
NAND2_X1 U_g3008C (.ZN(g3008C),.A2(g878C),.A1(g2444C));
NAND2_X1 U_I6836C (.ZN(I6836C),.A2(g806C),.A1(g3287C));
NAND2_X1 U_I5529C (.ZN(I5529C),.A2(I5528C),.A1(g1265C));
NAND2_X1 U_g10229C (.ZN(g10229C),.A2(I15609C),.A1(I15608C));
NAND2_X1 U_I13661C (.ZN(I13661C),.A2(I13659C),.A1(g8322C));
NAND2_X1 U_I13895C (.ZN(I13895C),.A2(I13893C),.A1(g1436C));
NAND2_X1 U_g2303C (.ZN(g2303C),.A2(I5343C),.A1(I5342C));
NAND2_X1 U_I12039C (.ZN(I12039C),.A2(I12038C),.A1(g5847C));
NAND2_X1 U_g5592C (.ZN(g5592C),.A2(I9008C),.A1(I9007C));
NAND2_X1 U_I12038C (.ZN(I12038C),.A2(g1466C),.A1(g5847C));
NAND2_X1 U_g3322C (.ZN(g3322C),.A2(I6489C),.A1(I6488C));
NAND2_X1 U_I8561C (.ZN(I8561C),.A2(g491C),.A1(g4227C));
NAND2_X1 U_I8527C (.ZN(I8527C),.A2(g481C),.A1(g4879C));
NAND2_X1 U_I12143C (.ZN(I12143C),.A2(g158C),.A1(g6000C));
NAND2_X1 U_I5619C (.ZN(I5619C),.A2(I5618C),.A1(g1766C));
NAND2_X1 U_g10386C (.ZN(g10386C),.A2(I15880C),.A1(I15879C));
NAND2_X1 U_I11980C (.ZN(I11980C),.A2(g1482C),.A1(g5820C));
NAND2_X1 U_I6837C (.ZN(I6837C),.A2(I6836C),.A1(g3287C));
NAND2_X1 U_I4973C (.ZN(I4973C),.A2(I4971C),.A1(g995C));
NAND2_X1 U_I13888C (.ZN(I13888C),.A2(I13886C),.A1(g1440C));
NAND2_X1 U_g7558C (.ZN(g7558C),.A2(I12004C),.A1(I12003C));
NAND2_X1 U_I17494C (.ZN(I17494C),.A2(I17492C),.A1(g3623C));
NAND2_X1 U_g11491C (.ZN(g11491C),.A2(I17494C),.A1(I17493C));
NAND2_X1 U_I16045C (.ZN(I16045C),.A2(I16044C),.A1(g833C));
NAND2_X1 U_I7684C (.ZN(I7684C),.A2(I7683C),.A1(g1023C));
NAND2_X1 U_g4130C (.ZN(g4130C),.A2(g2518C),.A1(FE_OFN352_g109C));
NAND2_X1 U_I8771C (.ZN(I8771C),.A2(I8770C),.A1(g4619C));
NAND2_X1 U_I13546C (.ZN(I13546C),.A2(I13544C),.A1(g8259C));
NAND2_X1 U_I13089C (.ZN(I13089C),.A2(g1840C),.A1(g8006C));
NAND2_X1 U_g2117C (.ZN(g2117C),.A2(I5025C),.A1(I5024C));
NAND2_X1 U_g5119C (.ZN(g5119C),.A2(I8515C),.A1(I8514C));
NAND2_X1 U_g5319C (.ZN(g5319C),.A2(I8805C),.A1(I8804C));
NAND2_X1 U_I15899C (.ZN(I15899C),.A2(I15898C),.A1(g857C));
NAND2_X1 U_I5606C (.ZN(I5606C),.A2(I5604C),.A1(g1153C));
NAND2_X1 U_I15898C (.ZN(I15898C),.A2(g10359C),.A1(g857C));
NAND2_X1 U_I16032C (.ZN(I16032C),.A2(I16030C),.A1(g10430C));
NAND2_X1 U_I17401C (.ZN(I17401C),.A2(I17400C),.A1(g11418C));
NAND2_X1 U_I13659C (.ZN(I13659C),.A2(g8322C),.A1(g1945C));
NAND2_X1 U_I8738C (.ZN(I8738C),.A2(g1121C),.A1(g4607C));
NAND2_X1 U_I13250C (.ZN(I13250C),.A2(I13248C),.A1(g8148C));
NAND2_X1 U_I15718C (.ZN(I15718C),.A2(I15716C),.A1(g10229C));
NAND2_X1 U_I9008C (.ZN(I9008C),.A2(I9006C),.A1(FE_OFN252_g1791C));
NAND2_X1 U_I6176C (.ZN(I6176C),.A2(g197C),.A1(g2177C));
NAND2_X1 U_I7865C (.ZN(I7865C),.A2(I7863C),.A1(g774C));
NAND2_X1 U_g5274C (.ZN(g5274C),.A2(I8730C),.A1(I8729C));
NAND2_X1 U_I5341C (.ZN(I5341C),.A2(g426C),.A1(g315C));
NAND2_X1 U_I17305C (.ZN(I17305C),.A2(g11231C),.A1(g11232C));
NAND2_X1 U_I17053C (.ZN(I17053C),.A2(I17051C),.A1(g11249C));
NAND2_X1 U_g5125C (.ZN(g5125C),.A2(I8529C),.A1(I8528C));
NAND2_X1 U_I12216C (.ZN(I12216C),.A2(I12214C),.A1(g2518C));
NAND2_X1 U_I6225C (.ZN(I6225C),.A2(I6224C),.A1(g2544C));
NAND2_X1 U_I5879C (.ZN(I5879C),.A2(I5878C),.A1(g2120C));
NAND2_X1 U_g3221C (.ZN(g3221C),.A2(g2564C),.A1(g1834C));
NAND2_X1 U_I14270C (.ZN(I14270C),.A2(g1822C),.A1(g8840C));
NAND2_X1 U_I6124C (.ZN(I6124C),.A2(g1419C),.A1(g2215C));
NAND2_X1 U_I6324C (.ZN(I6324C),.A2(I6322C),.A1(g1864C));
NAND2_X1 U_I13867C (.ZN(I13867C),.A2(g1403C),.A1(g8264C));
NAND2_X1 U_I13894C (.ZN(I13894C),.A2(I13893C),.A1(g8266C));
NAND2_X1 U_I6469C (.ZN(I6469C),.A2(I6467C),.A1(g2479C));
NAND2_X1 U_I8663C (.ZN(I8663C),.A2(I8662C),.A1(g4286C));
NAND2_X1 U_g7523C (.ZN(g7523C),.A2(I11909C),.A1(I11908C));
NAND2_X1 U_I6177C (.ZN(I6177C),.A2(I6176C),.A1(g2177C));
NAND2_X1 U_g5187C (.ZN(g5187C),.A2(I8591C),.A1(I8590C));
NAND2_X1 U_I6287C (.ZN(I6287C),.A2(g981C),.A1(g2091C));
NAND2_X1 U_I8762C (.ZN(I8762C),.A2(I8761C),.A1(g4616C));
NAND2_X1 U_I15871C (.ZN(I15871C),.A2(I15870C),.A1(g10291C));
NAND3_X1 U_g8840C (.ZN(g8840C),.A3(g8551C),.A2(g8541C),.A1(g8542C));
NAND2_X1 U_g2250C (.ZN(g2250C),.A2(I5265C),.A1(I5264C));
NAND2_X1 U_I8590C (.ZN(I8590C),.A2(I8589C),.A1(g4251C));
NAND2_X1 U_I6199C (.ZN(I6199C),.A2(g766C),.A1(g2525C));
NAND2_X1 U_I14218C (.ZN(I14218C),.A2(I14216C),.A1(g605C));
NAND2_X1 U_g8190C (.ZN(g8190C),.A2(g7978C),.A1(g6027C));
NAND2_X1 U_I5284C (.ZN(I5284C),.A2(I5282C),.A1(g762C));
NAND2_X1 U_I17485C (.ZN(I17485C),.A2(g11474C),.A1(g11233C));
NAND2_X1 U_I4965C (.ZN(I4965C),.A2(I4964C),.A1(g406C));
NAND2_X1 U_I5591C (.ZN(I5591C),.A2(g1703C),.A1(g1696C));
NAND2_X1 U_g8501C (.ZN(g8501C),.A2(g8366C),.A1(g3760C));
NAND2_X1 U_I15451C (.ZN(I15451C),.A2(g10019C),.A1(g10025C));
NAND2_X1 U_g8942C (.ZN(g8942C),.A2(FE_OFN200_g4921C),.A1(g8823C));
NAND2_X1 U_I13877C (.ZN(I13877C),.A2(I13876C),.A1(g8269C));
NAND2_X1 U_g7269C (.ZN(g7269C),.A2(I11510C),.A1(I11509C));
NAND2_X1 U_I4996C (.ZN(I4996C),.A2(I4995C),.A1(g416C));
NAND2_X1 U_I6144C (.ZN(I6144C),.A2(I6143C),.A1(g1976C));
NAND2_X1 U_I17567C (.ZN(I17567C),.A2(g1610C),.A1(g11496C));
NAND2_X1 U_g7572C (.ZN(g7572C),.A2(I12040C),.A1(I12039C));
NAND2_X1 U_I6207C (.ZN(I6207C),.A2(g802C),.A1(g5188C));
NAND2_X1 U_I14277C (.ZN(I14277C),.A2(g1828C),.A1(g8847C));
NAND2_X1 U_I16059C (.ZN(I16059C),.A2(I16058C),.A1(g841C));
NAND2_X1 U_I16025C (.ZN(I16025C),.A2(I16023C),.A1(FE_OFN253_g1786C));
NAND2_X1 U_I8563C (.ZN(I8563C),.A2(I8561C),.A1(g491C));
NAND2_X1 U_g3524C (.ZN(g3524C),.A2(g3221C),.A1(g3209C));
NAND2_X1 U_I16058C (.ZN(I16058C),.A2(g10441C),.A1(g841C));
NAND2_X1 U_I5204C (.ZN(I5204C),.A2(I5202C),.A1(g374C));
NAND2_X1 U_I6488C (.ZN(I6488C),.A2(I6487C),.A1(g2306C));
NAND4_X1 U_g3818C (.ZN(g3818C),.A4(g3003C),.A3(g2310C),.A2(g3071C),.A1(g3056C));
NAND2_X1 U_I16044C (.ZN(I16044C),.A2(g10432C),.A1(g833C));
NAND2_X1 U_g3717C (.ZN(g3717C),.A2(I6881C),.A1(I6880C));
NAND2_X1 U_I13077C (.ZN(I13077C),.A2(I13076C),.A1(g1872C));
NAND2_X1 U_g10043C (.ZN(g10043C),.A2(I15258C),.A1(I15257C));
NAND2_X1 U_I11280C (.ZN(I11280C),.A2(I11278C),.A1(g6485C));
NAND2_X1 U_I6825C (.ZN(I6825C),.A2(g770C),.A1(g3281C));
NAND2_X1 U_I4997C (.ZN(I4997C),.A2(I4995C),.A1(g309C));
NAND2_X1 U_I13300C (.ZN(I13300C),.A2(g8162C),.A1(g1936C));
NAND2_X1 U_I5323C (.ZN(I5323C),.A2(g1341C),.A1(g1336C));
NAND2_X1 U_I6136C (.ZN(I6136C),.A2(g378C),.A1(g2496C));
NAND2_X1 U_g5935C (.ZN(g5935C),.A2(I9559C),.A1(I9558C));
NAND2_X1 U_I5528C (.ZN(I5528C),.A2(g1015C),.A1(g1265C));
NAND2_X1 U_I6806C (.ZN(I6806C),.A2(I6805C),.A1(g3268C));
NAND2_X1 U_I5530C (.ZN(I5530C),.A2(I5528C),.A1(g1015C));
NAND2_X1 U_g10886C (.ZN(g10886C),.A2(g10805C),.A1(g10807C));
NAND2_X1 U_g3106C (.ZN(g3106C),.A2(I6324C),.A1(I6323C));
NAND2_X1 U_I13876C (.ZN(I13876C),.A2(g1444C),.A1(g8269C));
NAND2_X1 U_I6322C (.ZN(I6322C),.A2(g1864C),.A1(g2050C));
NAND2_X1 U_g3061C (.ZN(g3061C),.A2(g2374C),.A1(g611C));
NAND2_X1 U_g2439C (.ZN(g2439C),.A2(g1828C),.A1(g1814C));
NAND4_X1 U_g7947C (.ZN(g7947C),.A4(g7550C),.A3(FE_OFN91_g2172C),.A2(g7574C),.A1(g6941C));
NAND2_X1 U_I9576C (.ZN(I9576C),.A2(I9574C),.A1(g818C));
NAND2_X1 U_I13660C (.ZN(I13660C),.A2(I13659C),.A1(g1945C));
NAND2_X1 U_g3200C (.ZN(g3200C),.A2(g2061C),.A1(g1822C));
NAND2_X1 U_g4374C (.ZN(g4374C),.A2(I7685C),.A1(I7684C));
NAND2_X1 U_I11916C (.ZN(I11916C),.A2(I11914C),.A1(g1494C));
NAND2_X1 U_I5372C (.ZN(I5372C),.A2(I5371C),.A1(g971C));
NAND2_X1 U_g3003C (.ZN(g3003C),.A2(g2399C),.A1(g599C));
NAND2_X1 U_g8627C (.ZN(g8627C),.A2(I13888C),.A1(I13887C));
NAND2_X1 U_I5618C (.ZN(I5618C),.A2(FE_OFN247_g1771C),.A1(g1766C));
NAND2_X1 U_I6137C (.ZN(I6137C),.A2(I6136C),.A1(g2496C));
NAND2_X1 U_I5343C (.ZN(I5343C),.A2(I5341C),.A1(g426C));
NAND2_X1 U_I5282C (.ZN(I5282C),.A2(g762C),.A1(g758C));
NAND2_X1 U_I13307C (.ZN(I13307C),.A2(g617C),.A1(g8190C));
NAND2_X1 U_I13076C (.ZN(I13076C),.A2(g7963C),.A1(g1872C));
NAND2_X1 U_I6807C (.ZN(I6807C),.A2(I6805C),.A1(g471C));
NAND2_X1 U_I11243C (.ZN(I11243C),.A2(I11241C),.A1(g790C));
NAND2_X1 U_I17585C (.ZN(I17585C),.A2(I17584C),.A1(g11217C));
NAND2_X1 U_I12137C (.ZN(I12137C),.A2(I12136C),.A1(g6038C));
NAND2_X1 U_I7564C (.ZN(I7564C),.A2(I7562C),.A1(g654C));
NAND2_X1 U_g2970C (.ZN(g2970C),.A2(I6201C),.A1(I6200C));
NAND2_X1 U_g10144C (.ZN(g10144C),.A2(I15432C),.A1(I15431C));
NAND2_X1 U_I8788C (.ZN(I8788C),.A2(I8786C),.A1(g1141C));
NAND2_X1 U_g7054C (.ZN(g7054C),.A2(I11243C),.A1(I11242C));
NAND2_X1 U_I17052C (.ZN(I17052C),.A2(I17051C),.A1(g10923C));
NAND2_X1 U_g2120C (.ZN(g2120C),.A2(I5036C),.A1(I5035C));
NAND2_X1 U_g8616C (.ZN(g8616C),.A2(I13869C),.A1(I13868C));
NAND2_X1 U_I5202C (.ZN(I5202C),.A2(g374C),.A1(g369C));
NAND2_X1 U_I16088C (.ZN(I16088C),.A2(I16086C),.A1(g10430C));
NAND2_X1 U_I16024C (.ZN(I16024C),.A2(I16023C),.A1(g10438C));
NAND2_X1 U_g11490C (.ZN(g11490C),.A2(I17487C),.A1(I17486C));
NAND2_X1 U_I5518C (.ZN(I5518C),.A2(I5516C),.A1(g1019C));
NAND3_X1 U_g5118C (.ZN(g5118C),.A3(g4073C),.A2(g4806C),.A1(g2439C));
NAND2_X1 U_I12021C (.ZN(I12021C),.A2(I12019C),.A1(g166C));
NOR2_X1 U_g6392C (.ZN(g6392C),.A2(g5938C),.A1(g5859C));
NOR2_X1 U_g5938C (.ZN(g5938C),.A2(FE_OFN349_I6424C),.A1(g2273C));
NOR2_X1 U_g2478C (.ZN(g2478C),.A2(g1737C),.A1(g1610C));
NOR4_X1 U_g4278C (.ZN(g4278C),.A4(g3776C),.A3(FE_OFN254_g461C),.A2(FE_OFN248_g466C),.A1(g3800C));
NOR2_X1 U_g10383C (.ZN(g10383C),.A2(g3348C),.A1(I15514C));
NOR2_X1 U_g3118C (.ZN(g3118C),.A2(g2514C),.A1(g2521C));
NOR2_X1 U_g9815C (.ZN(g9815C),.A2(FE_OFN67_g9367C),.A1(FE_OFN68_g9392C));
NOR2_X1 U_g11077C (.ZN(g11077C),.A2(g10971C),.A1(g10970C));
NOR3_X1 U_g3879C (.ZN(g3879C),.A3(g2353C),.A2(g2354C),.A1(g3141C));
NOR2_X1 U_g10285C (.ZN(g10285C),.A2(FE_OFN350_g3121C),.A1(I15287C));
NOR2_X1 U_g11480C (.ZN(g11480C),.A2(g4567C),.A1(g11456C));
NOR2_X1 U_g4076C (.ZN(g4076C),.A2(I5254C),.A1(g1707C));
NOR2_X1 U_g10570C (.ZN(g10570C),.A2(g10324C),.A1(g10485C));
NOR2_X1 U_g10239C (.ZN(g10239C),.A2(I15287C),.A1(g9317C));
NOR2_X1 U_g10594C (.ZN(g10594C),.A2(g10521C),.A1(g10480C));
NOR2_X1 U_g9426C (.ZN(g9426C),.A2(FE_OFN50_g9030C),.A1(FE_OFN54_g9052C));
NOR2_X1 U_g10382C (.ZN(g10382C),.A2(g3348C),.A1(I15507C));
NOR4_X1 U_g4672C (.ZN(g4672C),.A4(g3479C),.A3(g1104C),.A2(g1107C),.A1(g3501C));
NOR2_X1 U_g5360C (.ZN(g5360C),.A2(FE_OFN308_I6424C),.A1(g105C));
NOR4_X1 U_g9387C (.ZN(g9387C),.A4(I14779C),.A3(g9223C),.A2(g9240C),.A1(g9010C));
NOR2_X1 U_g10438C (.ZN(g10438C),.A2(FE_OFN160_I6424C),.A1(I15500C));
NOR4_X1 U_g4613C (.ZN(g4613C),.A4(g1101C),.A3(g1104C),.A2(g3491C),.A1(FE_OFN240_g1110C));
NOR4_X1 U_g9391C (.ZN(g9391C),.A4(I14602C),.A3(FE_OFN39_g9223C),.A2(FE_OFN40_g9240C),.A1(g9010C));
NOR3_X1 U_g4572C (.ZN(g4572C),.A3(g3628C),.A2(g3408C),.A1(g3419C));
NOR3_X1 U_g9757C (.ZN(g9757C),.A3(FE_OFN72_g9292C),.A2(FE_OFN62_g9274C),.A1(FE_OFN32_g9454C));
NOR4_X1 U_g9874C (.ZN(g9874C),.A4(I15033C),.A3(g9579C),.A2(FE_OFN64_g9536C),.A1(g9519C));
NOR2_X1 U_g9654C (.ZN(g9654C),.A2(FE_OFN53_g9173C),.A1(FE_OFN46_g9125C));
NOR4_X1 U_g9880C (.ZN(g9880C),.A4(I15051C),.A3(g9579C),.A2(FE_OFN64_g9536C),.A1(g9751C));
NOR4_X1 U_g4873C (.ZN(g4873C),.A4(g3776C),.A3(FE_OFN254_g461C),.A2(FE_OFN248_g466C),.A1(FE_OFN250_g471C));
NOR2_X1 U_g2807C (.ZN(g2807C),.A2(g3629C),.A1(FE_OFN266_g18C));
NOR2_X1 U_g10441C (.ZN(g10441C),.A2(FE_OFN160_I6424C),.A1(I15510C));
NOR4_X1 U_g4639C (.ZN(g4639C),.A4(g1101C),.A3(g1104C),.A2(g1107C),.A1(g3501C));
NOR2_X1 U_g10435C (.ZN(g10435C),.A2(g3744C),.A1(I15510C));
NOR2_X1 U_g10849C (.ZN(g10849C),.A2(g2459C),.A1(g10739C));
NOR4_X1 U_g9606C (.ZN(g9606C),.A4(FE_OFN48_g9151C),.A3(FE_OFN52_g9173C),.A2(FE_OFN51_g9111C),.A1(FE_OFN45_g9125C));
NOR4_X1 U_g9879C (.ZN(g9879C),.A4(I15048C),.A3(g9563C),.A2(FE_OFN64_g9536C),.A1(g9747C));
NOR2_X1 U_g9506C (.ZN(g9506C),.A2(FE_OFN49_g9030C),.A1(FE_OFN56_g9052C));
NOR2_X1 U_g6155C (.ZN(g6155C),.A2(I5254C),.A1(g4974C));
NOR2_X1 U_g6355C (.ZN(g6355C),.A2(g6023C),.A1(g6032C));
NOR2_X1 U_g9591C (.ZN(g9591C),.A2(FE_OFN47_g9151C),.A1(FE_OFN44_g9125C));
NOR2_X1 U_g10359C (.ZN(g10359C),.A2(FE_OFN308_I6424C),.A1(I15290C));
NOR2_X1 U_g10434C (.ZN(g10434C),.A2(FE_OFN349_I6424C),.A1(I15514C));
NOR2_X1 U_g10291C (.ZN(g10291C),.A2(FE_OFN308_I6424C),.A1(I15287C));
NOR4_X1 U_g4227C (.ZN(g4227C),.A4(g2579C),.A3(FE_OFN254_g461C),.A2(g3793C),.A1(FE_OFN250_g471C));
NOR4_X1 U_g9667C (.ZN(g9667C),.A4(FE_OFN47_g9151C),.A3(FE_OFN52_g9173C),.A2(FE_OFN51_g9111C),.A1(FE_OFN45_g9125C));
NOR2_X1 U_g10563C (.ZN(g10563C),.A2(g10322C),.A1(g10484C));
NOR2_X1 U_g10324C (.ZN(g10324C),.A2(I15365C),.A1(g9317C));
NOR3_X1 U_g4455C (.ZN(g4455C),.A3(g3408C),.A2(g3419C),.A1(g3543C));
NOR4_X1 U_g9878C (.ZN(g9878C),.A4(I15045C),.A3(g9579C),.A2(FE_OFN64_g9536C),.A1(g9754C));
NOR2_X1 U_g10360C (.ZN(g10360C),.A2(FE_OFN350_g3121C),.A1(I15290C));
NOR4_X1 U_g9882C (.ZN(g9882C),.A4(I15057C),.A3(g9563C),.A2(FE_OFN64_g9536C),.A1(g9747C));
NOR4_X1 U_g4605C (.ZN(g4605C),.A4(g1101C),.A3(g3485C),.A2(g1107C),.A1(FE_OFN240_g1110C));
NOR2_X1 U_g10562C (.ZN(g10562C),.A2(g10529C),.A1(g10483C));
NOR2_X1 U_g5780C (.ZN(g5780C),.A2(FE_OFN200_g4921C),.A1(g3092C));
NOR2_X1 U_g10385C (.ZN(g10385C),.A2(g3348C),.A1(I15510C));
NOR4_X1 U_g4601C (.ZN(g4601C),.A4(g3479C),.A3(g1104C),.A2(g1107C),.A1(FE_OFN240_g1110C));
NOR2_X1 U_g5573C (.ZN(g5573C),.A2(g4432C),.A1(g4117C));
NOR2_X1 U_g5999C (.ZN(g5999C),.A2(FE_OFN349_I6424C),.A1(g2271C));
NOR3_X1 U_g9759C (.ZN(g9759C),.A3(FE_OFN71_g9292C),.A2(g9274C),.A1(g9454C));
NOR2_X1 U_g6037C (.ZN(g6037C),.A2(FE_OFN350_g3121C),.A1(g2297C));
NOR2_X1 U_g5034C (.ZN(g5034C),.A2(g3967C),.A1(g3524C));
NOR4_X1 U_g9881C (.ZN(g9881C),.A4(I15054C),.A3(g9579C),.A2(FE_OFN64_g9536C),.A1(g9516C));
NOR3_X1 U_g4276C (.ZN(g4276C),.A3(g2500C),.A2(g3261C),.A1(g4065C));
NOR4_X1 U_g4616C (.ZN(g4616C),.A4(g3479C),.A3(g1104C),.A2(g3491C),.A1(FE_OFN240_g1110C));
NOR2_X1 U_g10363C (.ZN(g10363C),.A2(FE_OFN308_I6424C),.A1(I15365C));
NOR2_X1 U_g2862C (.ZN(g2862C),.A2(g2305C),.A1(g2315C));
NOR3_X1 U_g9758C (.ZN(g9758C),.A3(FE_OFN71_g9292C),.A2(FE_OFN62_g9274C),.A1(FE_OFN32_g9454C));
NOR3_X1 U_g9589C (.ZN(g9589C),.A3(FE_OFN48_g9151C),.A2(FE_OFN52_g9173C),.A1(FE_OFN45_g9125C));
NOR2_X1 U_g9803C (.ZN(g9803C),.A2(g9367C),.A1(FE_OFN69_g9392C));
NOR2_X1 U_g10430C (.ZN(g10430C),.A2(FE_OFN349_I6424C),.A1(I15503C));
NOR2_X1 U_g10362C (.ZN(g10362C),.A2(g3744C),.A1(I15290C));
NOR2_X1 U_g2791C (.ZN(g2791C),.A2(g750C),.A1(g2187C));
NOR4_X1 U_g9605C (.ZN(g9605C),.A4(FE_OFN48_g9151C),.A3(FE_OFN52_g9173C),.A2(FE_OFN51_g9111C),.A1(FE_OFN46_g9125C));
NOR2_X1 U_g10436C (.ZN(g10436C),.A2(FE_OFN349_I6424C),.A1(I15510C));
NOR4_X1 U_g5556C (.ZN(g5556C),.A4(g2031C),.A3(g2299C),.A2(FE_OFN238_g1781C),.A1(g4787C));
NOR4_X1 U_g4286C (.ZN(g4286C),.A4(g2579C),.A3(g3784C),.A2(FE_OFN248_g466C),.A1(g3800C));
NOR2_X1 U_g4974C (.ZN(g4974C),.A2(g3714C),.A1(g4502C));
NOR2_X1 U_g9423C (.ZN(g9423C),.A2(FE_OFN49_g9030C),.A1(FE_OFN54_g9052C));
NOR2_X1 U_g5350C (.ZN(g5350C),.A2(FE_OFN160_I6424C),.A1(g3070C));
NOR4_X1 U_g2459C (.ZN(g2459C),.A4(g1648C),.A3(g1651C),.A2(g1642C),.A1(g1645C));
NOR2_X1 U_g10381C (.ZN(g10381C),.A2(g3348C),.A1(I15503C));
NOR4_X1 U_g4259C (.ZN(g4259C),.A4(g3776C),.A3(g3784C),.A2(g3793C),.A1(FE_OFN250_g471C));
NOR2_X1 U_g10522C (.ZN(g10522C),.A2(g10239C),.A1(g10401C));
NOR2_X1 U_g5392C (.ZN(g5392C),.A2(FE_OFN160_I6424C),.A1(g3086C));
NOR3_X1 U_g4122C (.ZN(g4122C),.A3(g2538C),.A2(g2410C),.A1(g3291C));
NOR2_X1 U_g6023C (.ZN(g6023C),.A2(FE_OFN160_I6424C),.A1(g2275C));
NOR2_X1 U_g3462C (.ZN(g3462C),.A2(g2795C),.A1(g2187C));
NOR4_X1 U_g4218C (.ZN(g4218C),.A4(g3776C),.A3(g3784C),.A2(FE_OFN248_g466C),.A1(FE_OFN250_g471C));
NOR4_X1 U_g4267C (.ZN(g4267C),.A4(g2579C),.A3(FE_OFN254_g461C),.A2(FE_OFN248_g466C),.A1(g3800C));
NOR4_X1 U_g4677C (.ZN(g4677C),.A4(g1101C),.A3(g3485C),.A2(g1107C),.A1(g3501C));
NOR2_X1 U_g9646C (.ZN(g9646C),.A2(FE_OFN47_g9151C),.A1(FE_OFN45_g9125C));
NOR2_X1 U_g2863C (.ZN(g2863C),.A2(g2309C),.A1(g2316C));
NOR2_X1 U_g6032C (.ZN(g6032C),.A2(FE_OFN349_I6424C),.A1(g3008C));
NOR4_X1 U_g9647C (.ZN(g9647C),.A4(FE_OFN48_g9151C),.A3(FE_OFN53_g9173C),.A2(FE_OFN51_g9111C),.A1(FE_OFN46_g9125C));
NOR2_X1 U_g5859C (.ZN(g5859C),.A2(FE_OFN349_I6424C),.A1(g2987C));
NOR2_X1 U_g10433C (.ZN(g10433C),.A2(g3744C),.A1(I15514C));
NOR4_X1 U_g4251C (.ZN(g4251C),.A4(g2579C),.A3(g3784C),.A2(g3793C),.A1(FE_OFN250_g471C));
NOR4_X1 U_g9876C (.ZN(g9876C),.A4(I15054C),.A3(FE_OFN56_g9052C),.A2(FE_OFN280_g9536C),.A1(g9522C));
NOR2_X1 U_g8303C (.ZN(g8303C),.A2(g4811C),.A1(g8209C));
NOR2_X1 U_g10429C (.ZN(g10429C),.A2(g3744C),.A1(I15503C));
NOR2_X1 U_g10428C (.ZN(g10428C),.A2(g3121C),.A1(I15503C));
NOR4_X1 U_g4234C (.ZN(g4234C),.A4(g3776C),.A3(FE_OFN254_g461C),.A2(g3793C),.A1(FE_OFN250_g471C));
NOR4_X1 U_g9877C (.ZN(g9877C),.A4(I15048C),.A3(g9569C),.A2(FE_OFN64_g9536C),.A1(g9512C));
NOR2_X1 U_g5186C (.ZN(g5186C),.A2(FE_OFN223_g4401C),.A1(g2047C));
NOR4_X1 U_g4619C (.ZN(g4619C),.A4(g1101C),.A3(g3485C),.A2(g3491C),.A1(FE_OFN240_g1110C));
NOR2_X1 U_g10432C (.ZN(g10432C),.A2(FE_OFN349_I6424C),.A1(I15507C));
NOR2_X1 U_g5345C (.ZN(g5345C),.A2(FE_OFN350_g3121C),.A1(g2067C));
NOR2_X1 U_g5763C (.ZN(g5763C),.A2(g5345C),.A1(g5350C));
NOR4_X1 U_g4879C (.ZN(g4879C),.A4(g2579C),.A3(g3784C),.A2(FE_OFN248_g466C),.A1(FE_OFN250_g471C));
NOR4_X1 U_g4607C (.ZN(g4607C),.A4(g3479C),.A3(g3485C),.A2(g1107C),.A1(FE_OFN240_g1110C));
NOR2_X1 U_g3107C (.ZN(g3107C),.A2(g2499C),.A1(g2501C));
NOR2_X1 U_g10322C (.ZN(g10322C),.A2(I15500C),.A1(g9317C));
NOR4_X1 U_g4630C (.ZN(g4630C),.A4(g3479C),.A3(g3485C),.A2(g3491C),.A1(FE_OFN240_g1110C));
NOR2_X1 U_g10364C (.ZN(g10364C),.A2(g3744C),.A1(I15507C));
SDFF_X1 U_g1289C (.Q(g1289C),.SE(test_seC),.SI(test_siC),.D(g4556C),.CK(CKC));
SDFF_X1 U_g1882C (.Q(g1882C),.SE(test_seC),.SI(g1289C),.D(g8943C),.CK(CKC));
SDFF_X1 U_g312C (.Q(g312C),.SE(test_seC),.SI(g1882C),.D(g255C),.CK(CKC));
SDFF_X1 U_g452C (.Q(g452C),.SE(test_seC),.SI(g312C),.D(g11257C),.CK(CKC));
SDFF_X1 U_g123C (.Q(g123C),.SE(test_seC),.SI(g452C),.D(g7032C),.CK(CKC));
SDFF_X1 U_g207C (.Q(g207C),.SE(test_seC),.SI(g123C),.D(g6830C),.CK(CKC));
SDFF_X1 U_g713C (.Q(g713C),.SE(test_seC),.SI(g207C),.D(g8920C),.CK(CKC));
SDFF_X1 U_g1153C (.Q(g1153C),.SE(test_seC),.SI(g713C),.D(g4340C),.CK(CKC));
SDFF_X1 U_g1209C (.Q(g1209C),.SE(test_seC),.SI(g1153C),.D(g10732C),.CK(CKC));
SDFF_X1 U_g1744C (.Q(g1744C),.SE(test_seC),.SI(g1209C),.D(g4239C),.CK(CKC));
SDFF_X1 U_g1558C (.Q(g1558C),.SE(test_seC),.SI(g1744C),.D(g6538C),.CK(CKC));
SDFF_X1 U_g695C (.Q(g695C),.SE(test_seC),.SI(g1558C),.D(g8887C),.CK(CKC));
SDFF_X1 U_g461C (.Q(g461C),.SE(test_seC),.SI(g695C),.D(g11372C),.CK(CKC));
SDFF_X1 U_g940C (.Q(g940C),.SE(test_seC),.SI(g461C),.D(g8260C),.CK(CKC));
SDFF_X1 U_g976C (.Q(g976C),.SE(test_seC),.SI(g940C),.D(g11391C),.CK(CKC));
SDFF_X1 U_g709C (.Q(g709C),.SE(test_seC),.SI(g976C),.D(g8432C),.CK(CKC));
SDFF_X1 U_g1092C (.Q(g1092C),.SE(test_seC),.SI(g709C),.D(g6088C),.CK(CKC));
SDFF_X1 U_g1574C (.Q(g1574C),.SE(test_seC),.SI(g1092C),.D(g6478C),.CK(CKC));
SDFF_X1 U_g1864C (.Q(g1864C),.SE(test_seC),.SI(g1574C),.D(g6795C),.CK(CKC));
SDFF_X1 U_g369C (.Q(g369C),.SE(test_seC),.SI(g1864C),.D(g11320C),.CK(CKC));
SDFF_X1 U_g1580C (.Q(g1580C),.SE(test_seC),.SI(g369C),.D(g6500C),.CK(CKC));
SDFF_X1 U_g1736C (.Q(g1736C),.SE(test_seC),.SI(g1580C),.D(g5392C),.CK(CKC));
SDFF_X1 U_g39C (.Q(g39C),.SE(test_seC),.SI(g1736C),.D(g10663C),.CK(CKC));
SDFF_X1 U_g1651C (.Q(g1651C),.SE(test_seC),.SI(g39C),.D(g10782C),.CK(CKC));
SDFF_X1 U_g1424C (.Q(g1424C),.SE(test_seC),.SI(g1651C),.D(g6216C),.CK(CKC));
SDFF_X1 U_g1737C (.Q(g1737C),.SE(test_seC),.SI(g1424C),.D(g1736C),.CK(CKC));
SDFF_X1 U_g1672C (.Q(g1672C),.SE(test_seC),.SI(g1737C),.D(g10858C),.CK(CKC));
SDFF_X1 U_g1077C (.Q(g1077C),.SE(test_seC),.SI(g1672C),.D(g5914C),.CK(CKC));
SDFF_X1 U_g1231C (.Q(g1231C),.SE(test_seC),.SI(g1077C),.D(g7590C),.CK(CKC));
SDFF_X1 U_g4C (.Q(g4C),.SE(test_seC),.SI(g1231C),.D(g6656C),.CK(CKC));
SDFF_X1 U_g774C (.Q(g774C),.SE(test_seC),.SI(g4C),.D(g6728C),.CK(CKC));
SDFF_X1 U_g1104C (.Q(g1104C),.SE(test_seC),.SI(g774C),.D(g5126C),.CK(CKC));
SDFF_X1 U_g1304C (.Q(g1304C),.SE(test_seC),.SI(g1104C),.D(g7290C),.CK(CKC));
SDFF_X1 U_g243C (.Q(g243C),.SE(test_seC),.SI(g1304C),.D(g6841C),.CK(CKC));
SDFF_X1 U_g1499C (.Q(g1499C),.SE(test_seC),.SI(g243C),.D(g8041C),.CK(CKC));
SDFF_X1 U_g1044C (.Q(g1044C),.SE(test_seC),.SI(g1499C),.D(g7106C),.CK(CKC));
SDFF_X1 U_g1444C (.Q(g1444C),.SE(test_seC),.SI(g1044C),.D(g8766C),.CK(CKC));
SDFF_X1 U_g757C (.Q(g757C),.SE(test_seC),.SI(g1444C),.D(g10788C),.CK(CKC));
SDFF_X1 U_g786C (.Q(g786C),.SE(test_seC),.SI(g757C),.D(g8019C),.CK(CKC));
SDFF_X1 U_g1543C (.Q(g1543C),.SE(test_seC),.SI(g786C),.D(g6545C),.CK(CKC));
SDFF_X1 U_g552C (.Q(g552C),.SE(test_seC),.SI(g1543C),.D(g10856C),.CK(CKC));
SDFF_X1 U_g315C (.Q(g315C),.SE(test_seC),.SI(g552C),.D(g256C),.CK(CKC));
SDFF_X1 U_g1534C (.Q(g1534C),.SE(test_seC),.SI(g315C),.D(g6533C),.CK(CKC));
SDFF_X1 U_g622C (.Q(g622C),.SE(test_seC),.SI(g1534C),.D(g8820C),.CK(CKC));
SDFF_X1 U_g1927C (.Q(g1927C),.SE(test_seC),.SI(g622C),.D(g8941C),.CK(CKC));
SDFF_X1 U_g1660C (.Q(g1660C),.SE(test_seC),.SI(g1927C),.D(g10859C),.CK(CKC));
SDFF_X1 U_g278C (.Q(g278C),.SE(test_seC),.SI(g1660C),.D(g6922C),.CK(CKC));
SDFF_X1 U_g1436C (.Q(g1436C),.SE(test_seC),.SI(g278C),.D(g8772C),.CK(CKC));
SDFF_X1 U_g718C (.Q(g718C),.SE(test_seC),.SI(g1436C),.D(g8433C),.CK(CKC));
SDFF_X1 U_g76C (.Q(g76C),.SE(test_seC),.SI(g718C),.D(g6526C),.CK(CKC));
SDFF_X1 U_g554C (.Q(g554C),.SE(test_seC),.SI(g76C),.D(g10793C),.CK(CKC));
SDFF_X1 U_g496C (.Q(g496C),.SE(test_seC),.SI(g554C),.D(g11333C),.CK(CKC));
SDFF_X1 U_g981C (.Q(g981C),.SE(test_seC),.SI(g496C),.D(g11392C),.CK(CKC));
SDFF_X1 U_g878C (.Q(g878C),.SE(test_seC),.SI(g981C),.D(g3506C),.CK(CKC));
SDFF_X1 U_g590C (.Q(g590C),.SE(test_seC),.SI(g878C),.D(g1713C),.CK(CKC));
SDFF_X1 U_g829C (.Q(g829C),.SE(test_seC),.SI(g590C),.D(g794C),.CK(CKC));
SDFF_X1 U_g1095C (.Q(g1095C),.SE(test_seC),.SI(g829C),.D(g6093C),.CK(CKC));
SDFF_X1 U_g704C (.Q(g704C),.SE(test_seC),.SI(g1095C),.D(g8889C),.CK(CKC));
SDFF_X1 U_g1265C (.Q(g1265C),.SE(test_seC),.SI(g704C),.D(g7302C),.CK(CKC));
SDFF_X1 U_g1786C (.Q(g1786C),.SE(test_seC),.SI(g1265C),.D(g6525C),.CK(CKC));
SDFF_X1 U_g682C (.Q(g682C),.SE(test_seC),.SI(g1786C),.D(g8429C),.CK(CKC));
SDFF_X1 U_g1296C (.Q(g1296C),.SE(test_seC),.SI(g682C),.D(g7292C),.CK(CKC));
SDFF_X1 U_g587C (.Q(g587C),.SE(test_seC),.SI(g1296C),.D(g104C),.CK(CKC));
SDFF_X1 U_g52C (.Q(g52C),.SE(test_seC),.SI(g587C),.D(g6621C),.CK(CKC));
SDFF_X1 U_g646C (.Q(g646C),.SE(test_seC),.SI(g52C),.D(g7134C),.CK(CKC));
SDFF_X1 U_g327C (.Q(g327C),.SE(test_seC),.SI(g646C),.D(g260C),.CK(CKC));
SDFF_X1 U_g1389C (.Q(g1389C),.SE(test_seC),.SI(g327C),.D(g6333C),.CK(CKC));
SDFF_X1 U_g1371C (.Q(g1371C),.SE(test_seC),.SI(g1389C),.D(g6826C),.CK(CKC));
SDFF_X1 U_g1956C (.Q(g1956C),.SE(test_seC),.SI(g1371C),.D(g1955C),.CK(CKC));
SDFF_X1 U_g1675C (.Q(g1675C),.SE(test_seC),.SI(g1956C),.D(g10860C),.CK(CKC));
SDFF_X1 U_g354C (.Q(g354C),.SE(test_seC),.SI(g1675C),.D(g11483C),.CK(CKC));
SDFF_X1 U_g113C (.Q(g113C),.SE(test_seC),.SI(g354C),.D(g6392C),.CK(CKC));
SDFF_X1 U_g639C (.Q(g639C),.SE(test_seC),.SI(g113C),.D(g7626C),.CK(CKC));
SDFF_X1 U_g1684C (.Q(g1684C),.SE(test_seC),.SI(g639C),.D(g10866C),.CK(CKC));
SDFF_X1 U_g1639C (.Q(g1639C),.SE(test_seC),.SI(g1684C),.D(g8193C),.CK(CKC));
SDFF_X1 U_g1791C (.Q(g1791C),.SE(test_seC),.SI(g1639C),.D(g6983C),.CK(CKC));
SDFF_X1 U_g248C (.Q(g248C),.SE(test_seC),.SI(g1791C),.D(g6839C),.CK(CKC));
SDFF_X1 U_g1707C (.Q(g1707C),.SE(test_seC),.SI(g248C),.D(g4076C),.CK(CKC));
SDFF_X1 U_g1759C (.Q(g1759C),.SE(test_seC),.SI(g1707C),.D(g4293C),.CK(CKC));
SDFF_X1 U_g351C (.Q(g351C),.SE(test_seC),.SI(g1759C),.D(g11482C),.CK(CKC));
SDFF_X1 U_g1957C (.Q(g1957C),.SE(test_seC),.SI(g351C),.D(g1956C),.CK(CKC));
SDFF_X1 U_g1604C (.Q(g1604C),.SE(test_seC),.SI(g1957C),.D(g6507C),.CK(CKC));
SDFF_X1 U_g1098C (.Q(g1098C),.SE(test_seC),.SI(g1604C),.D(g6096C),.CK(CKC));
SDFF_X1 U_g932C (.Q(g932C),.SE(test_seC),.SI(g1098C),.D(g8250C),.CK(CKC));
SDFF_X1 U_g126C (.Q(g126C),.SE(test_seC),.SI(g932C),.D(I8503C),.CK(CKC));
SDFF_X1 U_g1896C (.Q(g1896C),.SE(test_seC),.SI(g126C),.D(g8282C),.CK(CKC));
SDFF_X1 U_g736C (.Q(g736C),.SE(test_seC),.SI(g1896C),.D(g8435C),.CK(CKC));
SDFF_X1 U_g1019C (.Q(g1019C),.SE(test_seC),.SI(g736C),.D(g6924C),.CK(CKC));
SDFF_X1 U_g1362C (.Q(g1362C),.SE(test_seC),.SI(g1019C),.D(g6819C),.CK(CKC));
SDFF_X1 U_g745C (.Q(g745C),.SE(test_seC),.SI(g1362C),.D(g746C),.CK(CKC));
SDFF_X1 U_g1419C (.Q(g1419C),.SE(test_seC),.SI(g745C),.D(g6244C),.CK(CKC));
SDFF_X1 U_g58C (.Q(g58C),.SE(test_seC),.SI(g1419C),.D(g6627C),.CK(CKC));
SDFF_X1 U_g32C (.Q(g32C),.SE(test_seC),.SI(g58C),.D(g11286C),.CK(CKC));
SDFF_X1 U_g876C (.Q(g876C),.SE(test_seC),.SI(g32C),.D(g878C),.CK(CKC));
SDFF_X1 U_g1086C (.Q(g1086C),.SE(test_seC),.SI(g876C),.D(g6071C),.CK(CKC));
SDFF_X1 U_g1486C (.Q(g1486C),.SE(test_seC),.SI(g1086C),.D(g8046C),.CK(CKC));
SDFF_X1 U_g1730C (.Q(g1730C),.SE(test_seC),.SI(g1486C),.D(g10707C),.CK(CKC));
SDFF_X1 U_g1504C (.Q(g1504C),.SE(test_seC),.SI(g1730C),.D(g6198C),.CK(CKC));
SDFF_X1 U_g1470C (.Q(g1470C),.SE(test_seC),.SI(g1504C),.D(g8051C),.CK(CKC));
SDFF_X1 U_g822C (.Q(g822C),.SE(test_seC),.SI(g1470C),.D(g8024C),.CK(CKC));
SDFF_X1 U_g583C (.Q(g583C),.SE(test_seC),.SI(g822C),.D(g29C),.CK(CKC));
SDFF_X1 U_g1678C (.Q(g1678C),.SE(test_seC),.SI(g583C),.D(g10862C),.CK(CKC));
SDFF_X1 U_g174C (.Q(g174C),.SE(test_seC),.SI(g1678C),.D(g8050C),.CK(CKC));
SDFF_X1 U_g1766C (.Q(g1766C),.SE(test_seC),.SI(g174C),.D(g7133C),.CK(CKC));
SDFF_X1 U_g1801C (.Q(g1801C),.SE(test_seC),.SI(g1766C),.D(g7930C),.CK(CKC));
SDFF_X1 U_g186C (.Q(g186C),.SE(test_seC),.SI(g1801C),.D(g6832C),.CK(CKC));
SDFF_X1 U_g959C (.Q(g959C),.SE(test_seC),.SI(g186C),.D(g11308C),.CK(CKC));
SDFF_X1 U_g1169C (.Q(g1169C),.SE(test_seC),.SI(g959C),.D(g5189C),.CK(CKC));
SDFF_X1 U_g1007C (.Q(g1007C),.SE(test_seC),.SI(g1169C),.D(g6918C),.CK(CKC));
SDFF_X1 U_g1407C (.Q(g1407C),.SE(test_seC),.SI(g1007C),.D(g8769C),.CK(CKC));
SDFF_X1 U_g1059C (.Q(g1059C),.SE(test_seC),.SI(g1407C),.D(g7236C),.CK(CKC));
SDFF_X1 U_g1868C (.Q(g1868C),.SE(test_seC),.SI(g1059C),.D(g6909C),.CK(CKC));
SDFF_X1 U_g758C (.Q(g758C),.SE(test_seC),.SI(g1868C),.D(g4940C),.CK(CKC));
SDFF_X1 U_g1718C (.Q(g1718C),.SE(test_seC),.SI(g758C),.D(g5404C),.CK(CKC));
SDFF_X1 U_g396C (.Q(g396C),.SE(test_seC),.SI(g1718C),.D(g11265C),.CK(CKC));
SDFF_X1 U_g1015C (.Q(g1015C),.SE(test_seC),.SI(g396C),.D(g6930C),.CK(CKC));
SDFF_X1 U_g38C (.Q(g38C),.SE(test_seC),.SI(g1015C),.D(g10726C),.CK(CKC));
SDFF_X1 U_g632C (.Q(g632C),.SE(test_seC),.SI(g38C),.D(g4891C),.CK(CKC));
SDFF_X1 U_g1415C (.Q(g1415C),.SE(test_seC),.SI(g632C),.D(g6224C),.CK(CKC));
SDFF_X1 U_g1227C (.Q(g1227C),.SE(test_seC),.SI(g1415C),.D(g7586C),.CK(CKC));
SDFF_X1 U_g1721C (.Q(g1721C),.SE(test_seC),.SI(g1227C),.D(g10770C),.CK(CKC));
SDFF_X1 U_g882C (.Q(g882C),.SE(test_seC),.SI(g1721C),.D(g883C),.CK(CKC));
SDFF_X1 U_g16C (.Q(g16C),.SE(test_seC),.SI(g882C),.D(g3524C),.CK(CKC));
SDFF_X1 U_g284C (.Q(g284C),.SE(test_seC),.SI(g16C),.D(g6934C),.CK(CKC));
SDFF_X1 U_g426C (.Q(g426C),.SE(test_seC),.SI(g284C),.D(g11256C),.CK(CKC));
SDFF_X1 U_g219C (.Q(g219C),.SE(test_seC),.SI(g426C),.D(g6824C),.CK(CKC));
SDFF_X1 U_g1216C (.Q(g1216C),.SE(test_seC),.SI(g219C),.D(g1360C),.CK(CKC));
SDFF_X1 U_g806C (.Q(g806C),.SE(test_seC),.SI(g1216C),.D(g6126C),.CK(CKC));
SDFF_X1 U_g1428C (.Q(g1428C),.SE(test_seC),.SI(g806C),.D(g8767C),.CK(CKC));
SDFF_X1 U_g579C (.Q(g579C),.SE(test_seC),.SI(g1428C),.D(g102C),.CK(CKC));
SDFF_X1 U_g1564C (.Q(g1564C),.SE(test_seC),.SI(g579C),.D(g6546C),.CK(CKC));
SDFF_X1 U_g1741C (.Q(g1741C),.SE(test_seC),.SI(g1564C),.D(g4238C),.CK(CKC));
SDFF_X1 U_g225C (.Q(g225C),.SE(test_seC),.SI(g1741C),.D(g6823C),.CK(CKC));
SDFF_X1 U_g281C (.Q(g281C),.SE(test_seC),.SI(g225C),.D(g6928C),.CK(CKC));
SDFF_X1 U_g1308C (.Q(g1308C),.SE(test_seC),.SI(g281C),.D(g11602C),.CK(CKC));
SDFF_X1 U_g611C (.Q(g611C),.SE(test_seC),.SI(g1308C),.D(g9721C),.CK(CKC));
SDFF_X1 U_g631C (.Q(g631C),.SE(test_seC),.SI(g611C),.D(g4890C),.CK(CKC));
SDFF_X1 U_g1217C (.Q(g1217C),.SE(test_seC),.SI(g631C),.D(g9525C),.CK(CKC));
SDFF_X1 U_g1589C (.Q(g1589C),.SE(test_seC),.SI(g1217C),.D(g6524C),.CK(CKC));
SDFF_X1 U_g1466C (.Q(g1466C),.SE(test_seC),.SI(g1589C),.D(g8045C),.CK(CKC));
SDFF_X1 U_g1571C (.Q(g1571C),.SE(test_seC),.SI(g1466C),.D(g6469C),.CK(CKC));
SDFF_X1 U_g1861C (.Q(g1861C),.SE(test_seC),.SI(g1571C),.D(g6471C),.CK(CKC));
SDFF_X1 U_g1365C (.Q(g1365C),.SE(test_seC),.SI(g1861C),.D(g6821C),.CK(CKC));
SDFF_X1 U_g1448C (.Q(g1448C),.SE(test_seC),.SI(g1365C),.D(g11514C),.CK(CKC));
SDFF_X1 U_g1711C (.Q(g1711C),.SE(test_seC),.SI(g1448C),.D(g5403C),.CK(CKC));
SDFF_X1 U_g1133C (.Q(g1133C),.SE(test_seC),.SI(g1711C),.D(g4480C),.CK(CKC));
SDFF_X1 U_g1333C (.Q(g1333C),.SE(test_seC),.SI(g1133C),.D(g11610C),.CK(CKC));
SDFF_X1 U_g153C (.Q(g153C),.SE(test_seC),.SI(g1333C),.D(g7843C),.CK(CKC));
SDFF_X1 U_g962C (.Q(g962C),.SE(test_seC),.SI(g153C),.D(g11310C),.CK(CKC));
SDFF_X1 U_g766C (.Q(g766C),.SE(test_seC),.SI(g962C),.D(g5536C),.CK(CKC));
SDFF_X1 U_g588C (.Q(g588C),.SE(test_seC),.SI(g766C),.D(g28C),.CK(CKC));
SDFF_X1 U_g486C (.Q(g486C),.SE(test_seC),.SI(g588C),.D(g11331C),.CK(CKC));
SDFF_X1 U_g471C (.Q(g471C),.SE(test_seC),.SI(g486C),.D(g11380C),.CK(CKC));
SDFF_X1 U_g1397C (.Q(g1397C),.SE(test_seC),.SI(g471C),.D(g6838C),.CK(CKC));
SDFF_X1 U_g580C (.Q(g580C),.SE(test_seC),.SI(g1397C),.D(g103C),.CK(CKC));
SDFF_X1 U_g1950C (.Q(g1950C),.SE(test_seC),.SI(g580C),.D(g8288C),.CK(CKC));
SDFF_X1 U_g756C (.Q(g756C),.SE(test_seC),.SI(g1950C),.D(g755C),.CK(CKC));
SDFF_X1 U_g635C (.Q(g635C),.SE(test_seC),.SI(g756C),.D(g4892C),.CK(CKC));
SDFF_X1 U_g1101C (.Q(g1101C),.SE(test_seC),.SI(g635C),.D(g5390C),.CK(CKC));
SDFF_X1 U_g549C (.Q(g549C),.SE(test_seC),.SI(g1101C),.D(g10855C),.CK(CKC));
SDFF_X1 U_g1041C (.Q(g1041C),.SE(test_seC),.SI(g549C),.D(g7258C),.CK(CKC));
SDFF_X1 U_g105C (.Q(g105C),.SE(test_seC),.SI(g1041C),.D(g10898C),.CK(CKC));
SDFF_X1 U_g1669C (.Q(g1669C),.SE(test_seC),.SI(g105C),.D(g10865C),.CK(CKC));
SDFF_X1 U_g1368C (.Q(g1368C),.SE(test_seC),.SI(g1669C),.D(g6822C),.CK(CKC));
SDFF_X1 U_g1531C (.Q(g1531C),.SE(test_seC),.SI(g1368C),.D(g6528C),.CK(CKC));
SDFF_X1 U_g1458C (.Q(g1458C),.SE(test_seC),.SI(g1531C),.D(g6180C),.CK(CKC));
SDFF_X1 U_g572C (.Q(g572C),.SE(test_seC),.SI(g1458C),.D(g10718C),.CK(CKC));
SDFF_X1 U_g1011C (.Q(g1011C),.SE(test_seC),.SI(g572C),.D(g6912C),.CK(CKC));
SDFF_X1 U_g33C (.Q(g33C),.SE(test_seC),.SI(g1011C),.D(g10719C),.CK(CKC));
SDFF_X1 U_g1411C (.Q(g1411C),.SE(test_seC),.SI(g33C),.D(g6234C),.CK(CKC));
SDFF_X1 U_g1074C (.Q(g1074C),.SE(test_seC),.SI(g1411C),.D(g6099C),.CK(CKC));
SDFF_X1 U_g444C (.Q(g444C),.SE(test_seC),.SI(g1074C),.D(g11259C),.CK(CKC));
SDFF_X1 U_g1474C (.Q(g1474C),.SE(test_seC),.SI(g444C),.D(g8039C),.CK(CKC));
SDFF_X1 U_g1080C (.Q(g1080C),.SE(test_seC),.SI(g1474C),.D(g6059C),.CK(CKC));
SDFF_X1 U_g1713C (.Q(g1713C),.SE(test_seC),.SI(g1080C),.D(g5396C),.CK(CKC));
SDFF_X1 U_g333C (.Q(g333C),.SE(test_seC),.SI(g1713C),.D(g262C),.CK(CKC));
SDFF_X1 U_g269C (.Q(g269C),.SE(test_seC),.SI(g333C),.D(g6906C),.CK(CKC));
SDFF_X1 U_g401C (.Q(g401C),.SE(test_seC),.SI(g269C),.D(g11266C),.CK(CKC));
SDFF_X1 U_g1857C (.Q(g1857C),.SE(test_seC),.SI(g401C),.D(g11294C),.CK(CKC));
SDFF_X1 U_g9C (.Q(g9C),.SE(test_seC),.SI(g1857C),.D(g5421C),.CK(CKC));
SDFF_X1 U_g664C (.Q(g664C),.SE(test_seC),.SI(g9C),.D(g8649C),.CK(CKC));
SDFF_X1 U_g965C (.Q(g965C),.SE(test_seC),.SI(g664C),.D(g11312C),.CK(CKC));
SDFF_X1 U_g1400C (.Q(g1400C),.SE(test_seC),.SI(g965C),.D(g6840C),.CK(CKC));
SDFF_X1 U_g309C (.Q(g309C),.SE(test_seC),.SI(g1400C),.D(g254C),.CK(CKC));
SDFF_X1 U_g814C (.Q(g814C),.SE(test_seC),.SI(g309C),.D(g7202C),.CK(CKC));
SDFF_X1 U_g231C (.Q(g231C),.SE(test_seC),.SI(g814C),.D(g6834C),.CK(CKC));
SDFF_X1 U_g557C (.Q(g557C),.SE(test_seC),.SI(g231C),.D(g10795C),.CK(CKC));
SDFF_X1 U_g586C (.Q(g586C),.SE(test_seC),.SI(g557C),.D(g103C),.CK(CKC));
SDFF_X1 U_g869C (.Q(g869C),.SE(test_seC),.SI(g586C),.D(g875C),.CK(CKC));
SDFF_X1 U_g1383C (.Q(g1383C),.SE(test_seC),.SI(g869C),.D(g6831C),.CK(CKC));
SDFF_X1 U_g158C (.Q(g158C),.SE(test_seC),.SI(g1383C),.D(g8060C),.CK(CKC));
SDFF_X1 U_g627C (.Q(g627C),.SE(test_seC),.SI(g158C),.D(g4893C),.CK(CKC));
SDFF_X1 U_g1023C (.Q(g1023C),.SE(test_seC),.SI(g627C),.D(g7244C),.CK(CKC));
SDFF_X1 U_g259C (.Q(g259C),.SE(test_seC),.SI(g1023C),.D(g6026C),.CK(CKC));
SDFF_X1 U_g1361C (.Q(g1361C),.SE(test_seC),.SI(g259C),.D(g1206C),.CK(CKC));
SDFF_X1 U_g1327C (.Q(g1327C),.SE(test_seC),.SI(g1361C),.D(g11608C),.CK(CKC));
SDFF_X1 U_g654C (.Q(g654C),.SE(test_seC),.SI(g1327C),.D(g7660C),.CK(CKC));
SDFF_X1 U_g293C (.Q(g293C),.SE(test_seC),.SI(g654C),.D(g6911C),.CK(CKC));
SDFF_X1 U_g1346C (.Q(g1346C),.SE(test_seC),.SI(g293C),.D(g11640C),.CK(CKC));
SDFF_X1 U_g1633C (.Q(g1633C),.SE(test_seC),.SI(g1346C),.D(g8777C),.CK(CKC));
SDFF_X1 U_g1753C (.Q(g1753C),.SE(test_seC),.SI(g1633C),.D(g4274C),.CK(CKC));
SDFF_X1 U_g1508C (.Q(g1508C),.SE(test_seC),.SI(g1753C),.D(g6215C),.CK(CKC));
SDFF_X1 U_g1240C (.Q(g1240C),.SE(test_seC),.SI(g1508C),.D(g7297C),.CK(CKC));
SDFF_X1 U_g538C (.Q(g538C),.SE(test_seC),.SI(g1240C),.D(g11326C),.CK(CKC));
SDFF_X1 U_g416C (.Q(g416C),.SE(test_seC),.SI(g538C),.D(g11269C),.CK(CKC));
SDFF_X1 U_g542C (.Q(g542C),.SE(test_seC),.SI(g416C),.D(g11325C),.CK(CKC));
SDFF_X1 U_g1681C (.Q(g1681C),.SE(test_seC),.SI(g542C),.D(g10864C),.CK(CKC));
SDFF_X1 U_g374C (.Q(g374C),.SE(test_seC),.SI(g1681C),.D(g11290C),.CK(CKC));
SDFF_X1 U_g563C (.Q(g563C),.SE(test_seC),.SI(g374C),.D(g10798C),.CK(CKC));
SDFF_X1 U_g1914C (.Q(g1914C),.SE(test_seC),.SI(g563C),.D(g8284C),.CK(CKC));
SDFF_X1 U_g530C (.Q(g530C),.SE(test_seC),.SI(g1914C),.D(g11328C),.CK(CKC));
SDFF_X1 U_g575C (.Q(g575C),.SE(test_seC),.SI(g530C),.D(g10800C),.CK(CKC));
SDFF_X1 U_g1936C (.Q(g1936C),.SE(test_seC),.SI(g575C),.D(g8944C),.CK(CKC));
SDFF_X1 U_g55C (.Q(g55C),.SE(test_seC),.SI(g1936C),.D(g7183C),.CK(CKC));
SDFF_X1 U_g1117C (.Q(g1117C),.SE(test_seC),.SI(g55C),.D(g4465C),.CK(CKC));
SDFF_X1 U_g1317C (.Q(g1317C),.SE(test_seC),.SI(g1117C),.D(g1356C),.CK(CKC));
SDFF_X1 U_g357C (.Q(g357C),.SE(test_seC),.SI(g1317C),.D(g11484C),.CK(CKC));
SDFF_X1 U_g386C (.Q(g386C),.SE(test_seC),.SI(g357C),.D(g11263C),.CK(CKC));
SDFF_X1 U_g1601C (.Q(g1601C),.SE(test_seC),.SI(g386C),.D(g6501C),.CK(CKC));
SDFF_X1 U_g553C (.Q(g553C),.SE(test_seC),.SI(g1601C),.D(g10857C),.CK(CKC));
SDFF_X1 U_g166C (.Q(g166C),.SE(test_seC),.SI(g553C),.D(g6757C),.CK(CKC));
SDFF_X1 U_g501C (.Q(g501C),.SE(test_seC),.SI(g166C),.D(g11334C),.CK(CKC));
SDFF_X1 U_g262C (.Q(g262C),.SE(test_seC),.SI(g501C),.D(g6042C),.CK(CKC));
SDFF_X1 U_g1840C (.Q(g1840C),.SE(test_seC),.SI(g262C),.D(g8384C),.CK(CKC));
SDFF_X1 U_g70C (.Q(g70C),.SE(test_seC),.SI(g1840C),.D(g6653C),.CK(CKC));
SDFF_X1 U_g318C (.Q(g318C),.SE(test_seC),.SI(g70C),.D(g257C),.CK(CKC));
SDFF_X1 U_g1356C (.Q(g1356C),.SE(test_seC),.SI(g318C),.D(g5763C),.CK(CKC));
SDFF_X1 U_g794C (.Q(g794C),.SE(test_seC),.SI(g1356C),.D(g5849C),.CK(CKC));
SDFF_X1 U_g36C (.Q(g36C),.SE(test_seC),.SI(g794C),.D(g10722C),.CK(CKC));
SDFF_X1 U_g302C (.Q(g302C),.SE(test_seC),.SI(g36C),.D(g6929C),.CK(CKC));
SDFF_X1 U_g342C (.Q(g342C),.SE(test_seC),.SI(g302C),.D(g11488C),.CK(CKC));
SDFF_X1 U_g1250C (.Q(g1250C),.SE(test_seC),.SI(g342C),.D(g7299C),.CK(CKC));
SDFF_X1 U_g1163C (.Q(g1163C),.SE(test_seC),.SI(g1250C),.D(g4330C),.CK(CKC));
SDFF_X1 U_g1810C (.Q(g1810C),.SE(test_seC),.SI(g1163C),.D(g1958C),.CK(CKC));
SDFF_X1 U_g1032C (.Q(g1032C),.SE(test_seC),.SI(g1810C),.D(g7257C),.CK(CKC));
SDFF_X1 U_g1432C (.Q(g1432C),.SE(test_seC),.SI(g1032C),.D(g8775C),.CK(CKC));
SDFF_X1 U_g1053C (.Q(g1053C),.SE(test_seC),.SI(g1432C),.D(g7225C),.CK(CKC));
SDFF_X1 U_g1453C (.Q(g1453C),.SE(test_seC),.SI(g1053C),.D(g5770C),.CK(CKC));
SDFF_X1 U_g363C (.Q(g363C),.SE(test_seC),.SI(g1453C),.D(g11486C),.CK(CKC));
SDFF_X1 U_g330C (.Q(g330C),.SE(test_seC),.SI(g363C),.D(g261C),.CK(CKC));
SDFF_X1 U_g1157C (.Q(g1157C),.SE(test_seC),.SI(g330C),.D(g4338C),.CK(CKC));
SDFF_X1 U_g1357C (.Q(g1357C),.SE(test_seC),.SI(g1157C),.D(g4500C),.CK(CKC));
SDFF_X1 U_g35C (.Q(g35C),.SE(test_seC),.SI(g1357C),.D(g10721C),.CK(CKC));
SDFF_X1 U_g928C (.Q(g928C),.SE(test_seC),.SI(g35C),.D(g8147C),.CK(CKC));
SDFF_X1 U_g261C (.Q(g261C),.SE(test_seC),.SI(g928C),.D(g6038C),.CK(CKC));
SDFF_X1 U_g516C (.Q(g516C),.SE(test_seC),.SI(g261C),.D(g11337C),.CK(CKC));
SDFF_X1 U_g254C (.Q(g254C),.SE(test_seC),.SI(g516C),.D(g6045C),.CK(CKC));
SDFF_X1 U_g778C (.Q(g778C),.SE(test_seC),.SI(g254C),.D(g7191C),.CK(CKC));
SDFF_X1 U_g861C (.Q(g861C),.SE(test_seC),.SI(g778C),.D(g826C),.CK(CKC));
SDFF_X1 U_g1627C (.Q(g1627C),.SE(test_seC),.SI(g861C),.D(g8774C),.CK(CKC));
SDFF_X1 U_g1292C (.Q(g1292C),.SE(test_seC),.SI(g1627C),.D(g7293C),.CK(CKC));
SDFF_X1 U_g290C (.Q(g290C),.SE(test_seC),.SI(g1292C),.D(g6907C),.CK(CKC));
SDFF_X1 U_g1850C (.Q(g1850C),.SE(test_seC),.SI(g290C),.D(g4903C),.CK(CKC));
SDFF_X1 U_g770C (.Q(g770C),.SE(test_seC),.SI(g1850C),.D(g6123C),.CK(CKC));
SDFF_X1 U_g1583C (.Q(g1583C),.SE(test_seC),.SI(g770C),.D(g6506C),.CK(CKC));
SDFF_X1 U_g466C (.Q(g466C),.SE(test_seC),.SI(g1583C),.D(g11376C),.CK(CKC));
SDFF_X1 U_g1561C (.Q(g1561C),.SE(test_seC),.SI(g466C),.D(g6542C),.CK(CKC));
SDFF_X1 U_g1527C (.Q(g1527C),.SE(test_seC),.SI(g1561C),.D(I8503C),.CK(CKC));
SDFF_X1 U_g1546C (.Q(g1546C),.SE(test_seC),.SI(g1527C),.D(g6551C),.CK(CKC));
SDFF_X1 U_g287C (.Q(g287C),.SE(test_seC),.SI(g1546C),.D(g6901C),.CK(CKC));
SDFF_X1 U_g560C (.Q(g560C),.SE(test_seC),.SI(g287C),.D(g10797C),.CK(CKC));
SDFF_X1 U_g617C (.Q(g617C),.SE(test_seC),.SI(g560C),.D(g8505C),.CK(CKC));
SDFF_X1 U_g17C (.Q(g17C),.SE(test_seC),.SI(g617C),.D(g4117C),.CK(CKC));
SDFF_X1 U_g336C (.Q(g336C),.SE(test_seC),.SI(g17C),.D(g11647C),.CK(CKC));
SDFF_X1 U_g456C (.Q(g456C),.SE(test_seC),.SI(g336C),.D(g11340C),.CK(CKC));
SDFF_X1 U_g305C (.Q(g305C),.SE(test_seC),.SI(g456C),.D(g253C),.CK(CKC));
SDFF_X1 U_g345C (.Q(g345C),.SE(test_seC),.SI(g305C),.D(g11625C),.CK(CKC));
SDFF_X1 U_g8C (.Q(g8C),.SE(test_seC),.SI(g345C),.D(g636C),.CK(CKC));
SDFF_X1 U_g1771C (.Q(g1771C),.SE(test_seC),.SI(g8C),.D(g6502C),.CK(CKC));
SDFF_X1 U_g865C (.Q(g865C),.SE(test_seC),.SI(g1771C),.D(g7981C),.CK(CKC));
SDFF_X1 U_g255C (.Q(g255C),.SE(test_seC),.SI(g865C),.D(g6049C),.CK(CKC));
SDFF_X1 U_g1945C (.Q(g1945C),.SE(test_seC),.SI(g255C),.D(g8945C),.CK(CKC));
SDFF_X1 U_g1738C (.Q(g1738C),.SE(test_seC),.SI(g1945C),.D(g4231C),.CK(CKC));
SDFF_X1 U_g1478C (.Q(g1478C),.SE(test_seC),.SI(g1738C),.D(g8040C),.CK(CKC));
SDFF_X1 U_g1035C (.Q(g1035C),.SE(test_seC),.SI(g1478C),.D(g7203C),.CK(CKC));
SDFF_X1 U_g1959C (.Q(g1959C),.SE(test_seC),.SI(g1035C),.D(I5254C),.CK(CKC));
SDFF_X1 U_g1690C (.Q(g1690C),.SE(test_seC),.SI(g1959C),.D(g6155C),.CK(CKC));
SDFF_X1 U_g1482C (.Q(g1482C),.SE(test_seC),.SI(g1690C),.D(g8043C),.CK(CKC));
SDFF_X1 U_g1110C (.Q(g1110C),.SE(test_seC),.SI(g1482C),.D(g5173C),.CK(CKC));
SDFF_X1 U_g296C (.Q(g296C),.SE(test_seC),.SI(g1110C),.D(g6916C),.CK(CKC));
SDFF_X1 U_g1663C (.Q(g1663C),.SE(test_seC),.SI(g296C),.D(g10861C),.CK(CKC));
SDFF_X1 U_g700C (.Q(g700C),.SE(test_seC),.SI(g1663C),.D(g8431C),.CK(CKC));
SDFF_X1 U_g1762C (.Q(g1762C),.SE(test_seC),.SI(g700C),.D(g4309C),.CK(CKC));
SDFF_X1 U_g360C (.Q(g360C),.SE(test_seC),.SI(g1762C),.D(g11485C),.CK(CKC));
SDFF_X1 U_g192C (.Q(g192C),.SE(test_seC),.SI(g360C),.D(g6334C),.CK(CKC));
SDFF_X1 U_g1657C (.Q(g1657C),.SE(test_seC),.SI(g192C),.D(g10767C),.CK(CKC));
SDFF_X1 U_g722C (.Q(g722C),.SE(test_seC),.SI(g1657C),.D(g8923C),.CK(CKC));
SDFF_X1 U_g61C (.Q(g61C),.SE(test_seC),.SI(g722C),.D(g7189C),.CK(CKC));
SDFF_X1 U_g566C (.Q(g566C),.SE(test_seC),.SI(g61C),.D(g10799C),.CK(CKC));
SDFF_X1 U_g1394C (.Q(g1394C),.SE(test_seC),.SI(g566C),.D(g6747C),.CK(CKC));
SDFF_X1 U_g1089C (.Q(g1089C),.SE(test_seC),.SI(g1394C),.D(g6080C),.CK(CKC));
SDFF_X1 U_g883C (.Q(g883C),.SE(test_seC),.SI(g1089C),.D(g3381C),.CK(CKC));
SDFF_X1 U_g1071C (.Q(g1071C),.SE(test_seC),.SI(g883C),.D(g5910C),.CK(CKC));
SDFF_X1 U_g986C (.Q(g986C),.SE(test_seC),.SI(g1071C),.D(g11393C),.CK(CKC));
SDFF_X1 U_g971C (.Q(g971C),.SE(test_seC),.SI(g986C),.D(g11349C),.CK(CKC));
SDFF_X1 U_g1955C (.Q(g1955C),.SE(test_seC),.SI(g971C),.D(g83C),.CK(CKC));
SDFF_X1 U_g143C (.Q(g143C),.SE(test_seC),.SI(g1955C),.D(g6439C),.CK(CKC));
SDFF_X1 U_g1814C (.Q(g1814C),.SE(test_seC),.SI(g143C),.D(g9266C),.CK(CKC));
SDFF_X1 U_g1038C (.Q(g1038C),.SE(test_seC),.SI(g1814C),.D(g7245C),.CK(CKC));
SDFF_X1 U_g1212C (.Q(g1212C),.SE(test_seC),.SI(g1038C),.D(g1217C),.CK(CKC));
SDFF_X1 U_g1918C (.Q(g1918C),.SE(test_seC),.SI(g1212C),.D(g8940C),.CK(CKC));
SDFF_X1 U_g782C (.Q(g782C),.SE(test_seC),.SI(g1918C),.D(g7705C),.CK(CKC));
SDFF_X1 U_g1822C (.Q(g1822C),.SE(test_seC),.SI(g782C),.D(g9269C),.CK(CKC));
SDFF_X1 U_g237C (.Q(g237C),.SE(test_seC),.SI(g1822C),.D(g6820C),.CK(CKC));
SDFF_X1 U_g746C (.Q(g746C),.SE(test_seC),.SI(g237C),.D(g756C),.CK(CKC));
SDFF_X1 U_g1062C (.Q(g1062C),.SE(test_seC),.SI(g746C),.D(g7240C),.CK(CKC));
SDFF_X1 U_g1462C (.Q(g1462C),.SE(test_seC),.SI(g1062C),.D(g8042C),.CK(CKC));
SDFF_X1 U_g178C (.Q(g178C),.SE(test_seC),.SI(g1462C),.D(g6759C),.CK(CKC));
SDFF_X1 U_g366C (.Q(g366C),.SE(test_seC),.SI(g178C),.D(g11487C),.CK(CKC));
SDFF_X1 U_g837C (.Q(g837C),.SE(test_seC),.SI(g366C),.D(g802C),.CK(CKC));
SDFF_X1 U_g599C (.Q(g599C),.SE(test_seC),.SI(g837C),.D(g9124C),.CK(CKC));
SDFF_X1 U_g1854C (.Q(g1854C),.SE(test_seC),.SI(g599C),.D(g11293C),.CK(CKC));
SDFF_X1 U_g944C (.Q(g944C),.SE(test_seC),.SI(g1854C),.D(g11298C),.CK(CKC));
SDFF_X1 U_g1941C (.Q(g1941C),.SE(test_seC),.SI(g944C),.D(g8287C),.CK(CKC));
SDFF_X1 U_g170C (.Q(g170C),.SE(test_seC),.SI(g1941C),.D(g8047C),.CK(CKC));
SDFF_X1 U_g1520C (.Q(g1520C),.SE(test_seC),.SI(g170C),.D(g6205C),.CK(CKC));
SDFF_X1 U_g686C (.Q(g686C),.SE(test_seC),.SI(g1520C),.D(g8885C),.CK(CKC));
SDFF_X1 U_g953C (.Q(g953C),.SE(test_seC),.SI(g686C),.D(g11305C),.CK(CKC));
SDFF_X1 U_g1958C (.Q(g1958C),.SE(test_seC),.SI(g953C),.D(g5556C),.CK(CKC));
SDFF_X1 U_g40C (.Q(g40C),.SE(test_seC),.SI(g1958C),.D(g10664C),.CK(CKC));
SDFF_X1 U_g1765C (.Q(g1765C),.SE(test_seC),.SI(g40C),.D(g2478C),.CK(CKC));
SDFF_X1 U_g1733C (.Q(g1733C),.SE(test_seC),.SI(g1765C),.D(g10711C),.CK(CKC));
SDFF_X1 U_g1270C (.Q(g1270C),.SE(test_seC),.SI(g1733C),.D(g7303C),.CK(CKC));
SDFF_X1 U_g1610C (.Q(g1610C),.SE(test_seC),.SI(g1270C),.D(g5194C),.CK(CKC));
SDFF_X1 U_g1796C (.Q(g1796C),.SE(test_seC),.SI(g1610C),.D(g7541C),.CK(CKC));
SDFF_X1 U_g1324C (.Q(g1324C),.SE(test_seC),.SI(g1796C),.D(g11607C),.CK(CKC));
SDFF_X1 U_g1540C (.Q(g1540C),.SE(test_seC),.SI(g1324C),.D(g6541C),.CK(CKC));
SDFF_X1 U_g1377C (.Q(g1377C),.SE(test_seC),.SI(g1540C),.D(g6827C),.CK(CKC));
SDFF_X1 U_g1206C (.Q(g1206C),.SE(test_seC),.SI(g1377C),.D(g4114C),.CK(CKC));
SDFF_X1 U_g491C (.Q(g491C),.SE(test_seC),.SI(g1206C),.D(g11332C),.CK(CKC));
SDFF_X1 U_g1849C (.Q(g1849C),.SE(test_seC),.SI(g491C),.D(g4902C),.CK(CKC));
SDFF_X1 U_g213C (.Q(g213C),.SE(test_seC),.SI(g1849C),.D(g6828C),.CK(CKC));
SDFF_X1 U_g1781C (.Q(g1781C),.SE(test_seC),.SI(g213C),.D(g6516C),.CK(CKC));
SDFF_X1 U_g1900C (.Q(g1900C),.SE(test_seC),.SI(g1781C),.D(g8938C),.CK(CKC));
SDFF_X1 U_g1245C (.Q(g1245C),.SE(test_seC),.SI(g1900C),.D(g7298C),.CK(CKC));
SDFF_X1 U_g108C (.Q(g108C),.SE(test_seC),.SI(g1245C),.D(g11561C),.CK(CKC));
SDFF_X1 U_g630C (.Q(g630C),.SE(test_seC),.SI(g108C),.D(g6672C),.CK(CKC));
SDFF_X1 U_g148C (.Q(g148C),.SE(test_seC),.SI(g630C),.D(g8048C),.CK(CKC));
SDFF_X1 U_g833C (.Q(g833C),.SE(test_seC),.SI(g148C),.D(g798C),.CK(CKC));
SDFF_X1 U_g1923C (.Q(g1923C),.SE(test_seC),.SI(g833C),.D(g8285C),.CK(CKC));
SDFF_X1 U_g936C (.Q(g936C),.SE(test_seC),.SI(g1923C),.D(g8254C),.CK(CKC));
SDFF_X1 U_g1215C (.Q(g1215C),.SE(test_seC),.SI(g936C),.D(g5229C),.CK(CKC));
SDFF_X1 U_g1314C (.Q(g1314C),.SE(test_seC),.SI(g1215C),.D(g11604C),.CK(CKC));
SDFF_X1 U_g849C (.Q(g849C),.SE(test_seC),.SI(g1314C),.D(g814C),.CK(CKC));
SDFF_X1 U_g1336C (.Q(g1336C),.SE(test_seC),.SI(g849C),.D(g11636C),.CK(CKC));
SDFF_X1 U_g272C (.Q(g272C),.SE(test_seC),.SI(g1336C),.D(g6910C),.CK(CKC));
SDFF_X1 U_g1806C (.Q(g1806C),.SE(test_seC),.SI(g272C),.D(g8173C),.CK(CKC));
SDFF_X1 U_g826C (.Q(g826C),.SE(test_seC),.SI(g1806C),.D(g8245C),.CK(CKC));
SDFF_X1 U_g1065C (.Q(g1065C),.SE(test_seC),.SI(g826C),.D(g7242C),.CK(CKC));
SDFF_X1 U_g1887C (.Q(g1887C),.SE(test_seC),.SI(g1065C),.D(g8281C),.CK(CKC));
SDFF_X1 U_g37C (.Q(g37C),.SE(test_seC),.SI(g1887C),.D(g10724C),.CK(CKC));
SDFF_X1 U_g968C (.Q(g968C),.SE(test_seC),.SI(g37C),.D(g11314C),.CK(CKC));
SDFF_X1 U_g1845C (.Q(g1845C),.SE(test_seC),.SI(g968C),.D(g4905C),.CK(CKC));
SDFF_X1 U_g1137C (.Q(g1137C),.SE(test_seC),.SI(g1845C),.D(g4484C),.CK(CKC));
SDFF_X1 U_g1891C (.Q(g1891C),.SE(test_seC),.SI(g1137C),.D(g8937C),.CK(CKC));
SDFF_X1 U_g1255C (.Q(g1255C),.SE(test_seC),.SI(g1891C),.D(g7300C),.CK(CKC));
SDFF_X1 U_g257C (.Q(g257C),.SE(test_seC),.SI(g1255C),.D(g6002C),.CK(CKC));
SDFF_X1 U_g874C (.Q(g874C),.SE(test_seC),.SI(g257C),.D(g9507C),.CK(CKC));
SDFF_X1 U_g591C (.Q(g591C),.SE(test_seC),.SI(g874C),.D(g9110C),.CK(CKC));
SDFF_X1 U_g731C (.Q(g731C),.SE(test_seC),.SI(g591C),.D(g8926C),.CK(CKC));
SDFF_X1 U_g636C (.Q(g636C),.SE(test_seC),.SI(g731C),.D(g8631C),.CK(CKC));
SDFF_X1 U_g1218C (.Q(g1218C),.SE(test_seC),.SI(g636C),.D(g7632C),.CK(CKC));
SDFF_X1 U_g605C (.Q(g605C),.SE(test_seC),.SI(g1218C),.D(g9150C),.CK(CKC));
SDFF_X1 U_g79C (.Q(g79C),.SE(test_seC),.SI(g605C),.D(g6531C),.CK(CKC));
SDFF_X1 U_g182C (.Q(g182C),.SE(test_seC),.SI(g79C),.D(g6786C),.CK(CKC));
SDFF_X1 U_g950C (.Q(g950C),.SE(test_seC),.SI(g182C),.D(g11303C),.CK(CKC));
SDFF_X1 U_g1129C (.Q(g1129C),.SE(test_seC),.SI(g950C),.D(g4477C),.CK(CKC));
SDFF_X1 U_g857C (.Q(g857C),.SE(test_seC),.SI(g1129C),.D(g822C),.CK(CKC));
SDFF_X1 U_g448C (.Q(g448C),.SE(test_seC),.SI(g857C),.D(g11258C),.CK(CKC));
SDFF_X1 U_g1828C (.Q(g1828C),.SE(test_seC),.SI(g448C),.D(g9272C),.CK(CKC));
SDFF_X1 U_g1727C (.Q(g1727C),.SE(test_seC),.SI(g1828C),.D(g10773C),.CK(CKC));
SDFF_X1 U_g1592C (.Q(g1592C),.SE(test_seC),.SI(g1727C),.D(g6470C),.CK(CKC));
SDFF_X1 U_g1703C (.Q(g1703C),.SE(test_seC),.SI(g1592C),.D(g5083C),.CK(CKC));
SDFF_X1 U_g1932C (.Q(g1932C),.SE(test_seC),.SI(g1703C),.D(g8286C),.CK(CKC));
SDFF_X1 U_g1624C (.Q(g1624C),.SE(test_seC),.SI(g1932C),.D(g8773C),.CK(CKC));
SDFF_X1 U_g26C (.Q(g26C),.SE(test_seC),.SI(g1624C),.D(g4158C),.CK(CKC));
SDFF_X1 U_g1068C (.Q(g1068C),.SE(test_seC),.SI(g26C),.D(g6054C),.CK(CKC));
SDFF_X1 U_g578C (.Q(g578C),.SE(test_seC),.SI(g1068C),.D(g101C),.CK(CKC));
SDFF_X1 U_g440C (.Q(g440C),.SE(test_seC),.SI(g578C),.D(g11260C),.CK(CKC));
SDFF_X1 U_g476C (.Q(g476C),.SE(test_seC),.SI(g440C),.D(g11338C),.CK(CKC));
SDFF_X1 U_g119C (.Q(g119C),.SE(test_seC),.SI(g476C),.D(g5918C),.CK(CKC));
SDFF_X1 U_g668C (.Q(g668C),.SE(test_seC),.SI(g119C),.D(g8922C),.CK(CKC));
SDFF_X1 U_g139C (.Q(g139C),.SE(test_seC),.SI(g668C),.D(g8049C),.CK(CKC));
SDFF_X1 U_g1149C (.Q(g1149C),.SE(test_seC),.SI(g139C),.D(g4342C),.CK(CKC));
SDFF_X1 U_g34C (.Q(g34C),.SE(test_seC),.SI(g1149C),.D(g10720C),.CK(CKC));
SDFF_X1 U_g1848C (.Q(g1848C),.SE(test_seC),.SI(g34C),.D(g6755C),.CK(CKC));
SDFF_X1 U_g263C (.Q(g263C),.SE(test_seC),.SI(g1848C),.D(g6897C),.CK(CKC));
SDFF_X1 U_g818C (.Q(g818C),.SE(test_seC),.SI(g263C),.D(g7709C),.CK(CKC));
SDFF_X1 U_g1747C (.Q(g1747C),.SE(test_seC),.SI(g818C),.D(g4255C),.CK(CKC));
SDFF_X1 U_g802C (.Q(g802C),.SE(test_seC),.SI(g1747C),.D(g5543C),.CK(CKC));
SDFF_X1 U_g275C (.Q(g275C),.SE(test_seC),.SI(g802C),.D(g6915C),.CK(CKC));
SDFF_X1 U_g1524C (.Q(g1524C),.SE(test_seC),.SI(g275C),.D(g6513C),.CK(CKC));
SDFF_X1 U_g1577C (.Q(g1577C),.SE(test_seC),.SI(g1524C),.D(g6480C),.CK(CKC));
SDFF_X1 U_g810C (.Q(g810C),.SE(test_seC),.SI(g1577C),.D(g6733C),.CK(CKC));
SDFF_X1 U_g391C (.Q(g391C),.SE(test_seC),.SI(g810C),.D(g11264C),.CK(CKC));
SDFF_X1 U_g658C (.Q(g658C),.SE(test_seC),.SI(g391C),.D(g8973C),.CK(CKC));
SDFF_X1 U_g1386C (.Q(g1386C),.SE(test_seC),.SI(g658C),.D(g6833C),.CK(CKC));
SDFF_X1 U_g253C (.Q(g253C),.SE(test_seC),.SI(g1386C),.D(g5996C),.CK(CKC));
SDFF_X1 U_g875C (.Q(g875C),.SE(test_seC),.SI(g253C),.D(g9508C),.CK(CKC));
SDFF_X1 U_g1125C (.Q(g1125C),.SE(test_seC),.SI(g875C),.D(g4473C),.CK(CKC));
SDFF_X1 U_g201C (.Q(g201C),.SE(test_seC),.SI(g1125C),.D(g5755C),.CK(CKC));
SDFF_X1 U_g1280C (.Q(g1280C),.SE(test_seC),.SI(g201C),.D(g7295C),.CK(CKC));
SDFF_X1 U_g1083C (.Q(g1083C),.SE(test_seC),.SI(g1280C),.D(g6068C),.CK(CKC));
SDFF_X1 U_g650C (.Q(g650C),.SE(test_seC),.SI(g1083C),.D(g7137C),.CK(CKC));
SDFF_X1 U_g1636C (.Q(g1636C),.SE(test_seC),.SI(g650C),.D(g8779C),.CK(CKC));
SDFF_X1 U_g853C (.Q(g853C),.SE(test_seC),.SI(g1636C),.D(g818C),.CK(CKC));
SDFF_X1 U_g421C (.Q(g421C),.SE(test_seC),.SI(g853C),.D(g11270C),.CK(CKC));
SDFF_X1 U_g762C (.Q(g762C),.SE(test_seC),.SI(g421C),.D(g5529C),.CK(CKC));
SDFF_X1 U_g956C (.Q(g956C),.SE(test_seC),.SI(g762C),.D(g11306C),.CK(CKC));
SDFF_X1 U_g378C (.Q(g378C),.SE(test_seC),.SI(g956C),.D(g11291C),.CK(CKC));
SDFF_X1 U_g1756C (.Q(g1756C),.SE(test_seC),.SI(g378C),.D(g4283C),.CK(CKC));
SDFF_X1 U_g589C (.Q(g589C),.SE(test_seC),.SI(g1756C),.D(g29C),.CK(CKC));
SDFF_X1 U_g841C (.Q(g841C),.SE(test_seC),.SI(g589C),.D(g806C),.CK(CKC));
SDFF_X1 U_g1027C (.Q(g1027C),.SE(test_seC),.SI(g841C),.D(g6894C),.CK(CKC));
SDFF_X1 U_g1003C (.Q(g1003C),.SE(test_seC),.SI(g1027C),.D(g6902C),.CK(CKC));
SDFF_X1 U_g1403C (.Q(g1403C),.SE(test_seC),.SI(g1003C),.D(g8765C),.CK(CKC));
SDFF_X1 U_g1145C (.Q(g1145C),.SE(test_seC),.SI(g1403C),.D(g4498C),.CK(CKC));
SDFF_X1 U_g1107C (.Q(g1107C),.SE(test_seC),.SI(g1145C),.D(g5148C),.CK(CKC));
SDFF_X1 U_g1223C (.Q(g1223C),.SE(test_seC),.SI(g1107C),.D(g7581C),.CK(CKC));
SDFF_X1 U_g406C (.Q(g406C),.SE(test_seC),.SI(g1223C),.D(g11267C),.CK(CKC));
SDFF_X1 U_g1811C (.Q(g1811C),.SE(test_seC),.SI(g406C),.D(g10936C),.CK(CKC));
SDFF_X1 U_g1642C (.Q(g1642C),.SE(test_seC),.SI(g1811C),.D(g10784C),.CK(CKC));
SDFF_X1 U_g1047C (.Q(g1047C),.SE(test_seC),.SI(g1642C),.D(g7211C),.CK(CKC));
SDFF_X1 U_g1654C (.Q(g1654C),.SE(test_seC),.SI(g1047C),.D(g10765C),.CK(CKC));
SDFF_X1 U_g197C (.Q(g197C),.SE(test_seC),.SI(g1654C),.D(g6332C),.CK(CKC));
SDFF_X1 U_g1595C (.Q(g1595C),.SE(test_seC),.SI(g197C),.D(g6479C),.CK(CKC));
SDFF_X1 U_g1537C (.Q(g1537C),.SE(test_seC),.SI(g1595C),.D(g6537C),.CK(CKC));
SDFF_X1 U_g727C (.Q(g727C),.SE(test_seC),.SI(g1537C),.D(g8434C),.CK(CKC));
SDFF_X1 U_g999C (.Q(g999C),.SE(test_seC),.SI(g727C),.D(g6908C),.CK(CKC));
SDFF_X1 U_g798C (.Q(g798C),.SE(test_seC),.SI(g999C),.D(g6243C),.CK(CKC));
SDFF_X1 U_g481C (.Q(g481C),.SE(test_seC),.SI(g798C),.D(g11324C),.CK(CKC));
SDFF_X1 U_g754C (.Q(g754C),.SE(test_seC),.SI(g481C),.D(g3462C),.CK(CKC));
SDFF_X1 U_g1330C (.Q(g1330C),.SE(test_seC),.SI(g754C),.D(g11609C),.CK(CKC));
SDFF_X1 U_g845C (.Q(g845C),.SE(test_seC),.SI(g1330C),.D(g810C),.CK(CKC));
SDFF_X1 U_g790C (.Q(g790C),.SE(test_seC),.SI(g845C),.D(g8244C),.CK(CKC));
SDFF_X1 U_g1512C (.Q(g1512C),.SE(test_seC),.SI(g790C),.D(g8194C),.CK(CKC));
SDFF_X1 U_g114C (.Q(g114C),.SE(test_seC),.SI(g1512C),.D(g113C),.CK(CKC));
SDFF_X1 U_g1490C (.Q(g1490C),.SE(test_seC),.SI(g114C),.D(g8052C),.CK(CKC));
SDFF_X1 U_g1166C (.Q(g1166C),.SE(test_seC),.SI(g1490C),.D(g4325C),.CK(CKC));
SDFF_X1 U_g1056C (.Q(g1056C),.SE(test_seC),.SI(g1166C),.D(g7231C),.CK(CKC));
SDFF_X1 U_g348C (.Q(g348C),.SE(test_seC),.SI(g1056C),.D(g11481C),.CK(CKC));
SDFF_X1 U_g868C (.Q(g868C),.SE(test_seC),.SI(g348C),.D(g874C),.CK(CKC));
SDFF_X1 U_g1260C (.Q(g1260C),.SE(test_seC),.SI(g868C),.D(g7301C),.CK(CKC));
SDFF_X1 U_g260C (.Q(g260C),.SE(test_seC),.SI(g1260C),.D(g6035C),.CK(CKC));
SDFF_X1 U_g131C (.Q(g131C),.SE(test_seC),.SI(g260C),.D(g8059C),.CK(CKC));
SDFF_X1 U_g7C (.Q(g7C),.SE(test_seC),.SI(g131C),.D(g1854C),.CK(CKC));
SDFF_X1 U_g258C (.Q(g258C),.SE(test_seC),.SI(g7C),.D(g6015C),.CK(CKC));
SDFF_X1 U_g521C (.Q(g521C),.SE(test_seC),.SI(g258C),.D(g11330C),.CK(CKC));
SDFF_X1 U_g1318C (.Q(g1318C),.SE(test_seC),.SI(g521C),.D(g11605C),.CK(CKC));
SDFF_X1 U_g1872C (.Q(g1872C),.SE(test_seC),.SI(g1318C),.D(g8921C),.CK(CKC));
SDFF_X1 U_g677C (.Q(g677C),.SE(test_seC),.SI(g1872C),.D(g8883C),.CK(CKC));
SDFF_X1 U_g582C (.Q(g582C),.SE(test_seC),.SI(g677C),.D(g28C),.CK(CKC));
SDFF_X1 U_g1393C (.Q(g1393C),.SE(test_seC),.SI(g582C),.D(g6163C),.CK(CKC));
SDFF_X1 U_g1549C (.Q(g1549C),.SE(test_seC),.SI(g1393C),.D(g6523C),.CK(CKC));
SDFF_X1 U_g947C (.Q(g947C),.SE(test_seC),.SI(g1549C),.D(g11300C),.CK(CKC));
SDFF_X1 U_g1834C (.Q(g1834C),.SE(test_seC),.SI(g947C),.D(g9555C),.CK(CKC));
SDFF_X1 U_g1598C (.Q(g1598C),.SE(test_seC),.SI(g1834C),.D(g6481C),.CK(CKC));
SDFF_X1 U_g1121C (.Q(g1121C),.SE(test_seC),.SI(g1598C),.D(g4471C),.CK(CKC));
SDFF_X1 U_g1321C (.Q(g1321C),.SE(test_seC),.SI(g1121C),.D(g11606C),.CK(CKC));
SDFF_X1 U_g506C (.Q(g506C),.SE(test_seC),.SI(g1321C),.D(g11335C),.CK(CKC));
SDFF_X1 U_g546C (.Q(g546C),.SE(test_seC),.SI(g506C),.D(g10791C),.CK(CKC));
SDFF_X1 U_g1909C (.Q(g1909C),.SE(test_seC),.SI(g546C),.D(g8939C),.CK(CKC));
SDFF_X1 U_g755C (.Q(g755C),.SE(test_seC),.SI(g1909C),.D(g83C),.CK(CKC));
SDFF_X1 U_g1552C (.Q(g1552C),.SE(test_seC),.SI(g755C),.D(g6529C),.CK(CKC));
SDFF_X1 U_g584C (.Q(g584C),.SE(test_seC),.SI(g1552C),.D(g101C),.CK(CKC));
SDFF_X1 U_g1687C (.Q(g1687C),.SE(test_seC),.SI(g584C),.D(g10776C),.CK(CKC));
SDFF_X1 U_g1586C (.Q(g1586C),.SE(test_seC),.SI(g1687C),.D(g6514C),.CK(CKC));
SDFF_X1 U_g324C (.Q(g324C),.SE(test_seC),.SI(g1586C),.D(g259C),.CK(CKC));
SDFF_X1 U_g1141C (.Q(g1141C),.SE(test_seC),.SI(g324C),.D(g4490C),.CK(CKC));
SDFF_X1 U_g1570C (.Q(g1570C),.SE(test_seC),.SI(g1141C),.D(I8503C),.CK(CKC));
SDFF_X1 U_g1341C (.Q(g1341C),.SE(test_seC),.SI(g1570C),.D(g11639C),.CK(CKC));
SDFF_X1 U_g1710C (.Q(g1710C),.SE(test_seC),.SI(g1341C),.D(g4089C),.CK(CKC));
SDFF_X1 U_g1645C (.Q(g1645C),.SE(test_seC),.SI(g1710C),.D(g10785C),.CK(CKC));
SDFF_X1 U_g115C (.Q(g115C),.SE(test_seC),.SI(g1645C),.D(g6179C),.CK(CKC));
SDFF_X1 U_g135C (.Q(g135C),.SE(test_seC),.SI(g115C),.D(g8053C),.CK(CKC));
SDFF_X1 U_g525C (.Q(g525C),.SE(test_seC),.SI(g135C),.D(g11329C),.CK(CKC));
SDFF_X1 U_g581C (.Q(g581C),.SE(test_seC),.SI(g525C),.D(g104C),.CK(CKC));
SDFF_X1 U_g1607C (.Q(g1607C),.SE(test_seC),.SI(g581C),.D(g6515C),.CK(CKC));
SDFF_X1 U_g321C (.Q(g321C),.SE(test_seC),.SI(g1607C),.D(g258C),.CK(CKC));
SDFF_X1 U_g67C (.Q(g67C),.SE(test_seC),.SI(g321C),.D(g7204C),.CK(CKC));
SDFF_X1 U_g1275C (.Q(g1275C),.SE(test_seC),.SI(g67C),.D(g11443C),.CK(CKC));
SDFF_X1 U_g1311C (.Q(g1311C),.SE(test_seC),.SI(g1275C),.D(g11603C),.CK(CKC));
SDFF_X1 U_g1615C (.Q(g1615C),.SE(test_seC),.SI(g1311C),.D(g8770C),.CK(CKC));
SDFF_X1 U_g382C (.Q(g382C),.SE(test_seC),.SI(g1615C),.D(g11292C),.CK(CKC));
SDFF_X1 U_g1374C (.Q(g1374C),.SE(test_seC),.SI(g382C),.D(g6331C),.CK(CKC));
SDFF_X1 U_g266C (.Q(g266C),.SE(test_seC),.SI(g1374C),.D(g6900C),.CK(CKC));
SDFF_X1 U_g1284C (.Q(g1284C),.SE(test_seC),.SI(g266C),.D(g7294C),.CK(CKC));
SDFF_X1 U_g1380C (.Q(g1380C),.SE(test_seC),.SI(g1284C),.D(g6829C),.CK(CKC));
SDFF_X1 U_g673C (.Q(g673C),.SE(test_seC),.SI(g1380C),.D(g8428C),.CK(CKC));
SDFF_X1 U_g1853C (.Q(g1853C),.SE(test_seC),.SI(g673C),.D(g4904C),.CK(CKC));
SDFF_X1 U_g162C (.Q(g162C),.SE(test_seC),.SI(g1853C),.D(g8054C),.CK(CKC));
SDFF_X1 U_g411C (.Q(g411C),.SE(test_seC),.SI(g162C),.D(g11268C),.CK(CKC));
SDFF_X1 U_g431C (.Q(g431C),.SE(test_seC),.SI(g411C),.D(g11262C),.CK(CKC));
SDFF_X1 U_g1905C (.Q(g1905C),.SE(test_seC),.SI(g431C),.D(g8283C),.CK(CKC));
SDFF_X1 U_g1515C (.Q(g1515C),.SE(test_seC),.SI(g1905C),.D(g6193C),.CK(CKC));
SDFF_X1 U_g1630C (.Q(g1630C),.SE(test_seC),.SI(g1515C),.D(g8776C),.CK(CKC));
SDFF_X1 U_g49C (.Q(g49C),.SE(test_seC),.SI(g1630C),.D(g7143C),.CK(CKC));
SDFF_X1 U_g991C (.Q(g991C),.SE(test_seC),.SI(g49C),.D(g6898C),.CK(CKC));
SDFF_X1 U_g1300C (.Q(g1300C),.SE(test_seC),.SI(g991C),.D(g7291C),.CK(CKC));
SDFF_X1 U_g339C (.Q(g339C),.SE(test_seC),.SI(g1300C),.D(g11478C),.CK(CKC));
SDFF_X1 U_g256C (.Q(g256C),.SE(test_seC),.SI(g339C),.D(g6000C),.CK(CKC));
SDFF_X1 U_g1750C (.Q(g1750C),.SE(test_seC),.SI(g256C),.D(g4264C),.CK(CKC));
SDFF_X1 U_g585C (.Q(g585C),.SE(test_seC),.SI(g1750C),.D(g102C),.CK(CKC));
SDFF_X1 U_g1440C (.Q(g1440C),.SE(test_seC),.SI(g585C),.D(g8768C),.CK(CKC));
SDFF_X1 U_g1666C (.Q(g1666C),.SE(test_seC),.SI(g1440C),.D(g10863C),.CK(CKC));
SDFF_X1 U_g1528C (.Q(g1528C),.SE(test_seC),.SI(g1666C),.D(g6522C),.CK(CKC));
SDFF_X1 U_g1351C (.Q(g1351C),.SE(test_seC),.SI(g1528C),.D(g11641C),.CK(CKC));
SDFF_X1 U_g1648C (.Q(g1648C),.SE(test_seC),.SI(g1351C),.D(g10780C),.CK(CKC));
SDFF_X1 U_g127C (.Q(g127C),.SE(test_seC),.SI(g1648C),.D(g8044C),.CK(CKC));
SDFF_X1 U_g1618C (.Q(g1618C),.SE(test_seC),.SI(g127C),.D(g11579C),.CK(CKC));
SDFF_X1 U_g1235C (.Q(g1235C),.SE(test_seC),.SI(g1618C),.D(g7296C),.CK(CKC));
SDFF_X1 U_g299C (.Q(g299C),.SE(test_seC),.SI(g1235C),.D(g6923C),.CK(CKC));
SDFF_X1 U_g435C (.Q(g435C),.SE(test_seC),.SI(g299C),.D(g11261C),.CK(CKC));
SDFF_X1 U_g64C (.Q(g64C),.SE(test_seC),.SI(g435C),.D(g6638C),.CK(CKC));
SDFF_X1 U_g1555C (.Q(g1555C),.SE(test_seC),.SI(g64C),.D(g6534C),.CK(CKC));
SDFF_X1 U_g995C (.Q(g995C),.SE(test_seC),.SI(g1555C),.D(g6895C),.CK(CKC));
SDFF_X1 U_g1621C (.Q(g1621C),.SE(test_seC),.SI(g995C),.D(g8771C),.CK(CKC));
SDFF_X1 U_g1113C (.Q(g1113C),.SE(test_seC),.SI(g1621C),.D(g4506C),.CK(CKC));
SDFF_X1 U_g643C (.Q(g643C),.SE(test_seC),.SI(g1113C),.D(g7441C),.CK(CKC));
SDFF_X1 U_g1494C (.Q(g1494C),.SE(test_seC),.SI(g643C),.D(g8055C),.CK(CKC));
SDFF_X1 U_g1567C (.Q(g1567C),.SE(test_seC),.SI(g1494C),.D(g6468C),.CK(CKC));
SDFF_X1 U_g691C (.Q(g691C),.SE(test_seC),.SI(g1567C),.D(g8430C),.CK(CKC));
SDFF_X1 U_g534C (.Q(g534C),.SE(test_seC),.SI(g691C),.D(g11327C),.CK(CKC));
SDFF_X1 U_g1776C (.Q(g1776C),.SE(test_seC),.SI(g534C),.D(g6508C),.CK(CKC));
SDFF_X1 U_g569C (.Q(g569C),.SE(test_seC),.SI(g1776C),.D(g10717C),.CK(CKC));
SDFF_X1 U_g1160C (.Q(g1160C),.SE(test_seC),.SI(g569C),.D(g4334C),.CK(CKC));
SDFF_X1 U_g1360C (.Q(g1360C),.SE(test_seC),.SI(g1160C),.D(g9526C),.CK(CKC));
SDFF_X1 U_g1050C (.Q(g1050C),.SE(test_seC),.SI(g1360C),.D(g7218C),.CK(CKC));
SDFF_X1 U_g1C (.Q(g1C),.SE(test_seC),.SI(g1050C),.D(g6679C),.CK(CKC));
SDFF_X1 U_g511C (.Q(g511C),.SE(test_seC),.SI(g1C),.D(g11336C),.CK(CKC));
SDFF_X1 U_g1724C (.Q(g1724C),.SE(test_seC),.SI(g511C),.D(g10771C),.CK(CKC));
SDFF_X1 U_g12C (.Q(g12C),.SE(test_seC),.SI(g1724C),.D(g5445C),.CK(CKC));
SDFF_X1 U_g1878C (.Q(g1878C),.SE(test_seC),.SI(g12C),.D(g8559C),.CK(CKC));
SDFF_X1 U_g73C (.Q(g73C),.SE(test_seC),.SI(g1878C),.D(g7219C),.CK(CKC));
endmodule
